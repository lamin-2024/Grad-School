* File: Flip_Flop.pex.sp
* Created: Thu Nov 28 14:46:29 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.include "Flip_Flop.pex.sp.pex"
.subckt Flip_Flop  VSS Q VDD CLK D R
* 
* R	R
* D	D
* CLK	CLK
* VDD	VDD
* Q	Q
* VSS	VSS
XD0_noxref N_VSS_D0_noxref_pos N_VDD_D0_noxref_neg DIODENWX  AREA=4.61016e-11
+ PERIM=3.1764e-05
XMMN14 N_NET011_MMN14_d N_CLK_MMN14_g N_VSS_MMN14_s N_VSS_D0_noxref_pos NFET
+ L=6.2e-08 W=1.7e-06 AD=5.797e-13 AS=5.134e-13 PD=4.082e-06 PS=4.004e-06
+ NRD=0.0970588 NRS=0.0841176 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=3.02e-07 SB=3.41e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=0 PANW8=3.348e-15 PANW9=2.48e-14 PANW10=3.72e-14
XMMN13 N_NET07_MMN13_d N_NET011_MMN13_g N_VSS_MMN13_s N_VSS_D0_noxref_pos NFET
+ L=6.2e-08 W=1.7e-06 AD=4.114e-13 AS=8.262e-13 PD=3.884e-06 PS=4.372e-06
+ NRD=0.0782353 NRS=0.169412 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=4.86e-07 SB=2.42e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=0 PANW8=3.348e-15 PANW9=2.48e-14 PANW10=3.72e-14
XMMN3 NET5 N_D_MMN3_g N_VSS_MMN3_s N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=1.7e-06 AD=4.5305e-13 AS=5.1e-13 PD=2.233e-06 PS=4e-06 NRD=0.156765
+ NRS=0.0882353 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=3e-07
+ SB=3.394e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=3.348e-15 PANW9=2.48e-14 PANW10=3.72e-14
XMMN2 N_NET020_MMN2_d N_NET07_MMN2_g NET5 N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=1.7e-06 AD=2.55e-13 AS=4.5305e-13 PD=2e-06 PS=2.233e-06 NRD=0.0882353
+ NRS=0.156765 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=8.95e-07
+ SB=2.799e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=3.348e-15 PANW9=2.48e-14 PANW10=3.72e-14
XMMN5 N_NET020_MMN2_d N_NET011_MMN5_g NET054 N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=1.7e-06 AD=2.55e-13 AS=5.6695e-13 PD=2e-06 PS=2.367e-06 NRD=0.0882353
+ NRS=0.196176 M=1 NF=1 CNR_SWITCH=1 PCCRIT=0 PAR=1 PTWELL=0 SA=1.257e-06
+ SB=2.437e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=3.348e-15 PANW9=2.48e-14 PANW10=3.72e-14
XMMN4 NET054 N_NET027_MMN4_g N_VSS_MMN4_s N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=1.7e-06 AD=5.6695e-13 AS=4.2415e-13 PD=2.367e-06 PS=2.199e-06 NRD=0.196176
+ NRS=0.0876471 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.986e-06
+ SB=1.708e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=3.348e-15 PANW9=2.48e-14 PANW10=3.72e-14
XMMN0 N_NET027_MMN0_d N_NET020_MMN0_g N_VSS_MMN4_s N_VSS_D0_noxref_pos NFET
+ L=6.2e-08 W=1.7e-06 AD=4.2415e-13 AS=4.2415e-13 PD=2.199e-06 PS=2.199e-06
+ NRD=0.147059 NRS=0.205882 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=2.547e-06 SB=1.147e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=0 PANW8=3.348e-15 PANW9=2.48e-14 PANW10=3.72e-14
XMMN1 N_NET027_MMN0_d N_R_MMN1_g N_VSS_MMN1_s N_VSS_D0_noxref_pos NFET
+ L=6.2e-08 W=1.7e-06 AD=4.2415e-13 AS=9.962e-13 PD=2.199e-06 PS=4.572e-06
+ NRD=0.146471 NRS=0.237059 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=3.108e-06 SB=5.86e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=0 PANW8=3.348e-15 PANW9=2.48e-14 PANW10=3.72e-14
XMMN6 NET051 N_NET027_MMN6_g N_VSS_MMN6_s N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=1.7e-06 AD=3.944e-13 AS=5.78e-13 PD=2.164e-06 PS=4.08e-06 NRD=0.136471
+ NRS=0.0882353 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=3.4e-07
+ SB=3.001e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=3.348e-15 PANW9=2.48e-14 PANW10=3.72e-14
XMMN7 N_NET042_MMN7_d N_NET011_MMN7_g NET051 N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=1.7e-06 AD=2.55e-13 AS=3.944e-13 PD=2e-06 PS=2.164e-06 NRD=0.0882353
+ NRS=0.136471 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=8.66e-07
+ SB=2.475e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=3.348e-15 PANW9=2.48e-14 PANW10=3.72e-14
XMMN9 N_NET042_MMN7_d N_NET07_MMN9_g NET048 N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=1.7e-06 AD=2.55e-13 AS=6.052e-13 PD=2e-06 PS=2.412e-06 NRD=0.0882353
+ NRS=0.209412 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.228e-06
+ SB=2.113e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=3.348e-15 PANW9=2.48e-14 PANW10=3.72e-14
XMMN8 NET048 N_NET077_MMN8_g N_VSS_MMN8_s N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=1.7e-06 AD=6.052e-13 AS=3.3235e-13 PD=2.412e-06 PS=2.091e-06 NRD=0.209412
+ NRS=0.14 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=2.002e-06
+ SB=1.339e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=3.348e-15 PANW9=2.48e-14 PANW10=3.72e-14
XMMN10 N_NET077_MMN10_d N_NET042_MMN10_g N_VSS_MMN8_s N_VSS_D0_noxref_pos NFET
+ L=6.2e-08 W=1.7e-06 AD=4.2415e-13 AS=3.3235e-13 PD=2.199e-06 PS=2.091e-06
+ NRD=0.0882353 NRS=0.09 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=2.455e-06 SB=8.86e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=0 PANW8=3.348e-15 PANW9=2.48e-14 PANW10=3.72e-14
XMMN11 N_NET077_MMN10_d N_R_MMN11_g N_VSS_MMN11_s N_VSS_D0_noxref_pos NFET
+ L=6.2e-08 W=1.7e-06 AD=4.2415e-13 AS=5.525e-13 PD=2.199e-06 PS=4.05e-06
+ NRD=0.205294 NRS=0.0735294 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=3.016e-06 SB=3.25e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=0 PANW8=3.348e-15 PANW9=2.48e-14 PANW10=3.72e-14
XMMN12 N_Q_MMN12_d N_NET042_MMN12_g N_VSS_MMN12_s N_VSS_D0_noxref_pos NFET
+ L=6.2e-08 W=1.7e-06 AD=5.593e-13 AS=4.522e-13 PD=4.058e-06 PS=3.932e-06
+ NRD=0.131176 NRS=0.0794118 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=2.66e-07 SB=3.29e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=0 PANW8=3.348e-15 PANW9=2.48e-14 PANW10=3.72e-14
XMMP16 N_NET011_MMP16_d N_CLK_MMP16_g N_VDD_MMP16_s N_VDD_D0_noxref_neg PFET
+ L=6.2e-08 W=1.8e-06 AD=6.138e-13 AS=5.436e-13 PD=4.282e-06 PS=4.204e-06
+ NRD=0.09 NRS=0.0744444 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1
+ SA=3.02e-07 SB=3.41e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=1.13956e-13 PANW8=1.24e-14 PANW9=3.3418e-14 PANW10=7.44e-14
XMMP14 N_NET07_MMP14_d N_NET011_MMP14_g N_VDD_MMP14_s N_VDD_D0_noxref_neg PFET
+ L=6.2e-08 W=1.8e-06 AD=4.302e-13 AS=8.748e-13 PD=4.078e-06 PS=4.572e-06
+ NRD=0.0738889 NRS=0.168333 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1
+ SA=4.86e-07 SB=2.39e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=2.356e-15 PANW8=1.24e-14 PANW9=3.3418e-14 PANW10=1.86e-13
XMMP3 NET7 N_D_MMP3_g N_VDD_MMP3_s N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=1.8e-06 AD=4.797e-13 AS=5.4e-13 PD=2.333e-06 PS=4.2e-06 NRD=0.148056
+ NRS=0.0838889 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=3e-07
+ SB=3.394e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=2.356e-15 PANW8=1.24e-14 PANW9=3.3418e-14 PANW10=7.44e-14
XMMP2 N_NET020_MMP2_d N_NET011_MMP2_g NET7 N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=1.8e-06 AD=2.7e-13 AS=4.797e-13 PD=2.1e-06 PS=2.333e-06 NRD=0.0833333
+ NRS=0.148056 M=1 NF=1 CNR_SWITCH=1 PCCRIT=0 PAR=1 PTWELL=1 SA=8.95e-07
+ SB=2.799e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=2.356e-15 PANW8=1.24e-14 PANW9=3.3418e-14 PANW10=7.44e-14
XMMP5 N_NET020_MMP2_d N_NET07_MMP5_g NET053 N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=1.8e-06 AD=2.7e-13 AS=6.003e-13 PD=2.1e-06 PS=2.467e-06 NRD=0.0833333
+ NRS=0.185278 M=1 NF=1 CNR_SWITCH=1 PCCRIT=0 PAR=1 PTWELL=1 SA=1.257e-06
+ SB=2.437e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=2.356e-15 PANW8=1.24e-14 PANW9=3.3418e-14 PANW10=7.44e-14
XMMP6 NET053 N_NET027_MMP6_g N_VDD_MMP6_s N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=1.8e-06 AD=6.003e-13 AS=4.491e-13 PD=2.467e-06 PS=2.299e-06 NRD=0.185278
+ NRS=0.0822222 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.986e-06
+ SB=1.708e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=2.356e-15 PANW8=1.24e-14 PANW9=3.3418e-14 PANW10=7.44e-14
XMMP0 NET12 N_NET020_MMP0_g N_VDD_MMP6_s N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=1.8e-06 AD=4.491e-13 AS=4.491e-13 PD=2.299e-06 PS=2.299e-06 NRD=0.138611
+ NRS=0.195 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=2.547e-06
+ SB=1.147e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=2.356e-15 PANW8=1.24e-14 PANW9=3.3418e-14 PANW10=7.44e-14
XMMP1 N_NET027_MMP1_d N_R_MMP1_g NET12 N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=1.8e-06 AD=1.0548e-12 AS=4.491e-13 PD=4.772e-06 PS=2.299e-06 NRD=0.22
+ NRS=0.138611 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=3.108e-06
+ SB=5.86e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=2.356e-15 PANW8=1.24e-14 PANW9=3.3418e-14 PANW10=7.44e-14
XMMP7 NET052 N_NET027_MMP7_g N_VDD_MMP7_s N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=1.8e-06 AD=4.176e-13 AS=6.12e-13 PD=2.264e-06 PS=4.28e-06 NRD=0.128889
+ NRS=0.0838889 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=3.4e-07
+ SB=3.001e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=2.356e-15 PANW8=1.24e-14 PANW9=3.3418e-14 PANW10=7.44e-14
XMMP8 N_NET042_MMP8_d N_NET07_MMP8_g NET052 N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=1.8e-06 AD=2.7e-13 AS=4.176e-13 PD=2.1e-06 PS=2.264e-06 NRD=0.0833333
+ NRS=0.128889 M=1 NF=1 CNR_SWITCH=1 PCCRIT=0 PAR=1 PTWELL=1 SA=8.66e-07
+ SB=2.475e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=2.356e-15 PANW8=1.24e-14 PANW9=3.3418e-14 PANW10=7.44e-14
XMMP10 N_NET042_MMP8_d N_NET011_MMP10_g NET050 N_VDD_D0_noxref_neg PFET
+ L=6.2e-08 W=1.8e-06 AD=2.7e-13 AS=6.408e-13 PD=2.1e-06 PS=2.512e-06
+ NRD=0.0833333 NRS=0.197778 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1
+ SA=1.228e-06 SB=2.113e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=2.356e-15 PANW8=1.24e-14 PANW9=3.3418e-14 PANW10=7.44e-14
XMMP9 NET050 N_NET077_MMP9_g N_VDD_MMP9_s N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=1.8e-06 AD=6.408e-13 AS=3.519e-13 PD=2.512e-06 PS=2.191e-06 NRD=0.197778
+ NRS=0.132222 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=2.002e-06
+ SB=1.339e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=2.356e-15 PANW8=1.24e-14 PANW9=3.3418e-14 PANW10=7.44e-14
XMMP12 NET045 N_NET042_MMP12_g N_VDD_MMP9_s N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=1.8e-06 AD=4.491e-13 AS=3.519e-13 PD=2.299e-06 PS=2.191e-06 NRD=0.138611
+ NRS=0.085 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=2.455e-06
+ SB=8.86e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=2.356e-15 PANW8=1.24e-14 PANW9=3.3418e-14 PANW10=7.44e-14
XMMP11 N_NET077_MMP11_d N_R_MMP11_g NET045 N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=1.8e-06 AD=5.85e-13 AS=4.491e-13 PD=4.25e-06 PS=2.299e-06 NRD=0.103333
+ NRS=0.138611 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=3.016e-06
+ SB=3.25e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=2.356e-15 PANW8=1.24e-14 PANW9=3.3418e-14 PANW10=1.86e-13
XMMP13 N_Q_MMP13_d N_NET042_MMP13_g N_VDD_MMP13_s N_VDD_D0_noxref_neg PFET
+ L=6.2e-08 W=1.8e-06 AD=5.922e-13 AS=4.788e-13 PD=4.258e-06 PS=4.132e-06
+ NRD=0.123889 NRS=0.0688889 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1
+ SA=2.66e-07 SB=3.29e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=2.356e-15 PANW8=1.24e-13 PANW9=3.3418e-14 PANW10=7.44e-14
*
.include "Flip_Flop.pex.sp.FLIP_FLOP.pxi"
*
.ends
*
*
