* File: NOR2.pex.sp
* Created: Mon Dec  2 13:09:21 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.include "NOR2.pex.sp.pex"
.subckt NOR2  VSS OUT VDD A B
* 
* B	B
* A	A
* VDD	VDD
* OUT	OUT
* VSS	VSS
XD0_noxref N_VSS_D0_noxref_pos N_VDD_D0_noxref_neg DIODENWX  AREA=9.779e-12
+ PERIM=1.278e-05
XMMN0 N_OUT_MMN0_d N_A_MMN0_g N_VSS_MMN0_s N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=1.7e-06 AD=3.91e-13 AS=7.65e-13 PD=2.16e-06 PS=4.3e-06 NRD=0.139412
+ NRS=0.127059 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=4.5e-07
+ SB=1.29e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=3.348e-15 PANW9=2.48e-14 PANW10=3.72e-14
XMMN1 N_OUT_MMN0_d N_B_MMN1_g N_VSS_MMN1_s N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=1.7e-06 AD=3.91e-13 AS=1.3056e-12 PD=2.16e-06 PS=4.936e-06 NRD=0.131176
+ NRS=0.318824 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=9.72e-07
+ SB=7.68e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=3.348e-15 PANW9=2.48e-14 PANW10=3.72e-14
XMMP0 NET09 N_A_MMP0_g N_VDD_MMP0_s N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=1.8e-06 AD=4.14e-13 AS=8.1e-13 PD=2.26e-06 PS=4.5e-06 NRD=0.127778 NRS=0.125
+ M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=4.5e-07 SB=1.29e-06 SD=0
+ PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=2.356e-15 PANW8=1.24e-13
+ PANW9=3.1744e-14 PANW10=1.86e-13
XMMP1 N_OUT_MMP1_d N_B_MMP1_g NET09 N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=1.8e-06 AD=1.3824e-12 AS=4.14e-13 PD=5.136e-06 PS=2.26e-06 NRD=0.279444
+ NRS=0.127778 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=9.72e-07
+ SB=7.68e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=2.356e-15 PANW8=1.24e-14 PANW9=2.51344e-13 PANW10=7.8e-14
*
.include "NOR2.pex.sp.NOR2.pxi"
*
.ends
*
*
