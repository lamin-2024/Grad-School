* File: NOR3.pex.sp
* Created: Mon Dec  2 10:44:19 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.include "NOR3.pex.sp.pex"
.subckt NOR3  OUT VSS VDD A B C
* 
* C	C
* B	B
* A	A
* VDD	VDD
* VSS	VSS
* OUT	OUT
XD0_noxref N_VSS_D0_noxref_pos N_VDD_D0_noxref_neg DIODENWX  AREA=1.17925e-11
+ PERIM=1.3826e-05
XMMN0 N_OUT_MMN0_d N_A_MMN0_g N_VSS_MMN0_s N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=1.7e-06 AD=7.65e-13 AS=3.91e-13 PD=4.3e-06 PS=2.16e-06 NRD=0.127059
+ NRS=0.138824 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=4.5e-07
+ SB=1.813e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=3.348e-15 PANW9=2.48e-14 PANW10=3.72e-14
XMMN1 N_OUT_MMN1_d N_B_MMN1_g N_VSS_MMN0_s N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=1.7e-06 AD=3.893e-13 AS=3.91e-13 PD=2.158e-06 PS=2.16e-06 NRD=0.131765
+ NRS=0.131765 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=9.72e-07
+ SB=1.291e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=3.348e-15 PANW9=2.48e-14 PANW10=3.72e-14
XMMN2 N_OUT_MMN1_d N_C_MMN2_g N_VSS_MMN2_s N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=1.7e-06 AD=3.893e-13 AS=1.3107e-12 PD=2.158e-06 PS=4.942e-06 NRD=0.137647
+ NRS=0.244706 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.492e-06
+ SB=7.71e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=3.348e-15 PANW9=2.48e-14 PANW10=3.72e-14
XMMP4 NET012 N_A_MMP4_g N_VDD_MMP4_s N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=1.8e-06 AD=4.14e-13 AS=8.1e-13 PD=2.26e-06 PS=4.5e-06 NRD=0.127778 NRS=0.125
+ M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=4.5e-07 SB=1.813e-06 SD=0
+ PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=2.356e-15 PANW8=1.24e-13
+ PANW9=3.1744e-14 PANW10=7.44e-14
XMMP0 NET09 N_B_MMP0_g NET012 N_VDD_D0_noxref_neg PFET L=6.2e-08 W=1.8e-06
+ AD=4.122e-13 AS=4.14e-13 PD=2.258e-06 PS=2.26e-06 NRD=0.127222 NRS=0.127778
+ M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=9.72e-07 SB=1.291e-06 SD=0
+ PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=2.356e-15 PANW8=1.24e-14
+ PANW9=1.39744e-13 PANW10=1.896e-13
XMMP1 N_OUT_MMP1_d N_C_MMP1_g NET09 N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=1.8e-06 AD=1.3878e-12 AS=4.122e-13 PD=5.142e-06 PS=2.258e-06 NRD=0.215556
+ NRS=0.127222 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.492e-06
+ SB=7.71e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=2.356e-15 PANW8=1.24e-14 PANW9=1.43344e-13 PANW10=1.86e-13
*
.include "NOR3.pex.sp.NOR3.pxi"
*
.ends
*
*
