module INV(IN, OUT);
input IN;
output OUT;
//assign OUT = ~IN;
endmodule

module NAND2(A, B, OUT);
input A, B;
output OUT;
//assign OUT = ~(A & B);
endmodule

module NAND3(A, B, C, OUT);
input A, B, C;
output OUT;
//assign OUT = ~(A & B & C);
endmodule

module NAND4(A, B, C, D, OUT);
input A, B, C, D;
output OUT;
//assign OUT = ~(A & B & C & D);
endmodule

module NOR2(A, B, OUT);
input A, B;
output OUT;
//assign OUT = ~(A | B);
endmodule

module NOR3(A, B, C, OUT);
input A, B, C;
output OUT;
//assign OUT = ~(A | B | C);
endmodule

module XOR2(A, B, OUT);
input A, B;
output OUT;
//assign OUT = (A ^ B);
endmodule

module AOI12(A, B, C, OUT);
input A, B, C;
output OUT;
//assign OUT = ~(A | (B & C));
endmodule

module AOI22(A, B, C, D, OUT);
input A, B, C, D;
output OUT;
//assign OUT = ~((A & B) | (C & D));
endmodule

module OAI12(A, B, C, OUT);
input A, B, C;
output OUT;
//assign OUT = ~(A & (B | C));
endmodule

module OAI22(A, B, C, D, OUT);
input A, B, C, D;
output OUT;
//assign OUT = ~((A | B) & (C | D));
endmodule

module Flip_Flop( D, CLK, R, Q);
input D, CLK, R;
output Q;
reg Q;
/*always @(posedge gclk or negedge rnot)
  if (rnot == 1'b0)
    Q = 1'b0;
  else
    Q = D;*/
endmodule



/////////////////////////////////////////////////////////////
// Created by: Synopsys DC Expert(TM) in wire load mode
// Version   : O-2018.06-SP1
// Date      : Mon Dec  2 15:14:46 2024
/////////////////////////////////////////////////////////////


module FIR_Filter_Project1_1 ( Data_out, Data_in, clock, reset );
  output [19:0] Data_out;
  input [7:0] Data_in;
  input clock, reset;
  wire   \Samples[13][7] , \Samples[13][6] , \Samples[13][5] ,
         \Samples[13][4] , \Samples[13][3] , \Samples[13][2] ,
         \Samples[13][1] , \Samples[13][0] , \Samples[12][7] ,
         \Samples[12][6] , \Samples[12][5] , \Samples[12][4] ,
         \Samples[12][3] , \Samples[12][2] , \Samples[12][1] ,
         \Samples[12][0] , \Samples[11][7] , \Samples[11][6] ,
         \Samples[11][5] , \Samples[11][4] , \Samples[11][3] ,
         \Samples[11][2] , \Samples[11][1] , \Samples[11][0] ,
         \Samples[10][7] , \Samples[10][6] , \Samples[10][5] ,
         \Samples[10][4] , \Samples[10][3] , \Samples[10][2] ,
         \Samples[10][1] , \Samples[10][0] , \Samples[9][7] , \Samples[9][6] ,
         \Samples[9][5] , \Samples[9][4] , \Samples[9][3] , \Samples[9][2] ,
         \Samples[9][1] , \Samples[9][0] , \Samples[8][7] , \Samples[8][6] ,
         \Samples[8][5] , \Samples[8][4] , \Samples[8][3] , \Samples[8][2] ,
         \Samples[8][1] , \Samples[8][0] , \Samples[7][7] , \Samples[7][6] ,
         \Samples[7][5] , \Samples[7][4] , \Samples[7][3] , \Samples[7][2] ,
         \Samples[7][1] , \Samples[7][0] , \Samples[6][7] , \Samples[6][6] ,
         \Samples[6][5] , \Samples[6][4] , \Samples[6][3] , \Samples[6][2] ,
         \Samples[6][1] , \Samples[6][0] , \Samples[5][7] , \Samples[5][6] ,
         \Samples[5][5] , \Samples[5][4] , \Samples[5][3] , \Samples[5][2] ,
         \Samples[5][1] , \Samples[5][0] , \Samples[4][7] , \Samples[4][6] ,
         \Samples[4][5] , \Samples[4][4] , \Samples[4][3] , \Samples[4][2] ,
         \Samples[4][1] , \Samples[4][0] , \Samples[3][7] , \Samples[3][6] ,
         \Samples[3][5] , \Samples[3][4] , \Samples[3][3] , \Samples[3][2] ,
         \Samples[3][1] , \Samples[3][0] , \Samples[2][7] , \Samples[2][6] ,
         \Samples[2][5] , \Samples[2][4] , \Samples[2][3] , \Samples[2][2] ,
         \Samples[2][1] , \Samples[2][0] , \Samples[1][7] , \Samples[1][6] ,
         \Samples[1][5] , \Samples[1][4] , \Samples[1][3] , \Samples[1][2] ,
         \Samples[1][1] , \Samples[1][0] , \Samples[0][7] , \Samples[0][6] ,
         \Samples[0][5] , \Samples[0][4] , \Samples[0][3] , \Samples[0][2] ,
         \Samples[0][1] , \Samples[0][0] , N3, N4, N5, N6, N7, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40,
         N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54,
         N55, N56, N57, N58, N59, N60, N63, N64, N65, N66, N67, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, \PR_mul[14][9] ,
         \PR_mul[14][8] , \PR_mul[14][7] , \PR_mul[14][6] , \PR_mul[14][5] ,
         \PR_mul[14][4] , \PR_mul[14][3] , \PR_mul[14][2] , \PR_mul[13][11] ,
         \PR_mul[13][10] , \PR_mul[13][9] , \PR_mul[13][8] , \PR_mul[13][7] ,
         \PR_mul[13][6] , \PR_mul[13][5] , \PR_mul[13][4] , \PR_mul[13][3] ,
         \PR_mul[13][2] , \PR_mul[12][11] , \PR_mul[12][10] , \PR_mul[12][9] ,
         \PR_mul[12][8] , \PR_mul[12][7] , \PR_mul[12][6] , \PR_mul[12][5] ,
         \PR_mul[12][4] , \PR_mul[12][3] , \PR_mul[12][2] , \PR_mul[12][1] ,
         \PR_mul[12][0] , \PR_mul[11][10] , \PR_mul[11][9] , \PR_mul[11][8] ,
         \PR_mul[11][7] , \PR_mul[11][6] , \PR_mul[11][5] , \PR_mul[11][4] ,
         \PR_mul[11][3] , \PR_mul[10][10] , \PR_mul[10][9] , \PR_mul[10][8] ,
         \PR_mul[10][7] , \PR_mul[10][6] , \PR_mul[10][5] , \PR_mul[10][4] ,
         \PR_mul[10][3] , \PR_mul[10][2] , \PR_mul[10][1] , \PR_mul[10][0] ,
         \PR_mul[9][9] , \PR_mul[9][8] , \PR_mul[9][7] , \PR_mul[9][6] ,
         \PR_mul[9][5] , \PR_mul[9][4] , \PR_mul[9][3] , \PR_mul[9][2] ,
         \PR_mul[8][11] , \PR_mul[8][10] , \PR_mul[8][9] , \PR_mul[8][8] ,
         \PR_mul[8][7] , \PR_mul[8][6] , \PR_mul[8][5] , \PR_mul[8][4] ,
         \PR_mul[8][3] , \PR_mul[8][2] , \PR_mul[7][11] , \PR_mul[7][10] ,
         \PR_mul[7][9] , \PR_mul[7][8] , \PR_mul[7][7] , \PR_mul[7][6] ,
         \PR_mul[7][5] , \PR_mul[7][4] , \PR_mul[7][3] , \PR_mul[7][2] ,
         \PR_mul[7][1] , \PR_mul[7][0] , \PR_mul[6][10] , \PR_mul[6][9] ,
         \PR_mul[6][8] , \PR_mul[6][7] , \PR_mul[6][6] , \PR_mul[6][5] ,
         \PR_mul[6][4] , \PR_mul[6][3] , \PR_mul[5][10] , \PR_mul[5][9] ,
         \PR_mul[5][8] , \PR_mul[5][7] , \PR_mul[5][6] , \PR_mul[5][5] ,
         \PR_mul[5][4] , \PR_mul[5][3] , \PR_mul[5][2] , \PR_mul[5][1] ,
         \PR_mul[5][0] , \PR_mul[4][9] , \PR_mul[4][8] , \PR_mul[4][7] ,
         \PR_mul[4][6] , \PR_mul[4][5] , \PR_mul[4][4] , \PR_mul[4][3] ,
         \PR_mul[4][2] , \PR_mul[3][11] , \PR_mul[3][10] , \PR_mul[3][9] ,
         \PR_mul[3][8] , \PR_mul[3][7] , \PR_mul[3][6] , \PR_mul[3][5] ,
         \PR_mul[3][4] , \PR_mul[3][3] , \PR_mul[3][2] , \PR_mul[2][11] ,
         \PR_mul[2][10] , \PR_mul[2][9] , \PR_mul[2][8] , \PR_mul[2][7] ,
         \PR_mul[2][6] , \PR_mul[2][5] , \PR_mul[2][4] , \PR_mul[2][3] ,
         \PR_mul[2][2] , \PR_mul[2][1] , \PR_mul[2][0] , \PR_mul[1][10] ,
         \PR_mul[1][9] , \PR_mul[1][8] , \PR_mul[1][7] , \PR_mul[1][6] ,
         \PR_mul[1][5] , \PR_mul[1][4] , \PR_mul[1][3] , \PR_mul[0][10] ,
         \PR_mul[0][9] , \PR_mul[0][8] , \PR_mul[0][7] , \PR_mul[0][6] ,
         \PR_mul[0][5] , \PR_mul[0][4] , \PR_mul[0][3] , N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119,
         \PR_add[13][19] , \PR_add[13][18] , \PR_add[13][17] ,
         \PR_add[13][16] , \PR_add[13][15] , \PR_add[13][14] ,
         \PR_add[13][13] , \PR_add[13][12] , \PR_add[13][11] ,
         \PR_add[13][10] , \PR_add[13][9] , \PR_add[13][8] , \PR_add[13][7] ,
         \PR_add[13][6] , \PR_add[13][5] , \PR_add[13][4] , \PR_add[13][3] ,
         \PR_add[13][2] , \PR_add[13][1] , \PR_add[13][0] , \PR_add[12][19] ,
         \PR_add[12][18] , \PR_add[12][17] , \PR_add[12][16] ,
         \PR_add[12][15] , \PR_add[12][14] , \PR_add[12][13] ,
         \PR_add[12][12] , \PR_add[12][11] , \PR_add[12][10] , \PR_add[12][9] ,
         \PR_add[12][8] , \PR_add[12][7] , \PR_add[12][6] , \PR_add[12][5] ,
         \PR_add[12][4] , \PR_add[12][3] , \PR_add[12][2] , \PR_add[11][19] ,
         \PR_add[11][18] , \PR_add[11][17] , \PR_add[11][16] ,
         \PR_add[11][15] , \PR_add[11][14] , \PR_add[11][13] ,
         \PR_add[11][12] , \PR_add[11][11] , \PR_add[11][10] , \PR_add[11][9] ,
         \PR_add[11][8] , \PR_add[11][7] , \PR_add[11][6] , \PR_add[11][5] ,
         \PR_add[11][4] , \PR_add[11][3] , \PR_add[11][2] , \PR_add[11][1] ,
         \PR_add[10][19] , \PR_add[10][18] , \PR_add[10][17] ,
         \PR_add[10][16] , \PR_add[10][15] , \PR_add[10][14] ,
         \PR_add[10][13] , \PR_add[10][12] , \PR_add[10][11] ,
         \PR_add[10][10] , \PR_add[10][9] , \PR_add[10][8] , \PR_add[10][7] ,
         \PR_add[10][6] , \PR_add[10][5] , \PR_add[10][4] , \PR_add[10][3] ,
         \PR_add[10][2] , \PR_add[10][1] , \PR_add[10][0] , \PR_add[9][19] ,
         \PR_add[9][18] , \PR_add[9][17] , \PR_add[9][16] , \PR_add[9][15] ,
         \PR_add[9][14] , \PR_add[9][13] , \PR_add[9][12] , \PR_add[9][11] ,
         \PR_add[9][10] , \PR_add[9][9] , \PR_add[9][8] , \PR_add[9][7] ,
         \PR_add[9][6] , \PR_add[9][5] , \PR_add[9][4] , \PR_add[9][3] ,
         \PR_add[8][19] , \PR_add[8][18] , \PR_add[8][17] , \PR_add[8][16] ,
         \PR_add[8][15] , \PR_add[8][14] , \PR_add[8][13] , \PR_add[8][12] ,
         \PR_add[8][11] , \PR_add[8][10] , \PR_add[8][9] , \PR_add[8][8] ,
         \PR_add[8][7] , \PR_add[8][6] , \PR_add[8][5] , \PR_add[8][4] ,
         \PR_add[8][3] , \PR_add[8][2] , \PR_add[8][1] , \PR_add[8][0] ,
         \PR_add[7][19] , \PR_add[7][18] , \PR_add[7][17] , \PR_add[7][16] ,
         \PR_add[7][15] , \PR_add[7][14] , \PR_add[7][13] , \PR_add[7][12] ,
         \PR_add[7][11] , \PR_add[7][10] , \PR_add[7][9] , \PR_add[7][8] ,
         \PR_add[7][7] , \PR_add[7][6] , \PR_add[7][5] , \PR_add[7][4] ,
         \PR_add[7][3] , \PR_add[7][2] , \PR_add[6][19] , \PR_add[6][18] ,
         \PR_add[6][17] , \PR_add[6][16] , \PR_add[6][15] , \PR_add[6][14] ,
         \PR_add[6][13] , \PR_add[6][12] , \PR_add[6][11] , \PR_add[6][10] ,
         \PR_add[6][9] , \PR_add[6][8] , \PR_add[6][7] , \PR_add[6][6] ,
         \PR_add[6][5] , \PR_add[6][4] , \PR_add[6][3] , \PR_add[6][2] ,
         \PR_add[6][1] , \PR_add[5][19] , \PR_add[5][18] , \PR_add[5][17] ,
         \PR_add[5][16] , \PR_add[5][15] , \PR_add[5][14] , \PR_add[5][13] ,
         \PR_add[5][12] , \PR_add[5][11] , \PR_add[5][10] , \PR_add[5][9] ,
         \PR_add[5][8] , \PR_add[5][7] , \PR_add[5][6] , \PR_add[5][5] ,
         \PR_add[5][4] , \PR_add[5][3] , \PR_add[5][2] , \PR_add[5][1] ,
         \PR_add[5][0] , \PR_add[4][19] , \PR_add[4][18] , \PR_add[4][17] ,
         \PR_add[4][16] , \PR_add[4][15] , \PR_add[4][14] , \PR_add[4][13] ,
         \PR_add[4][12] , \PR_add[4][11] , \PR_add[4][10] , \PR_add[4][9] ,
         \PR_add[4][8] , \PR_add[4][7] , \PR_add[4][6] , \PR_add[4][5] ,
         \PR_add[4][4] , \PR_add[4][3] , \PR_add[3][19] , \PR_add[3][18] ,
         \PR_add[3][17] , \PR_add[3][16] , \PR_add[3][15] , \PR_add[3][14] ,
         \PR_add[3][13] , \PR_add[3][12] , \PR_add[3][11] , \PR_add[3][10] ,
         \PR_add[3][9] , \PR_add[3][8] , \PR_add[3][7] , \PR_add[3][6] ,
         \PR_add[3][5] , \PR_add[3][4] , \PR_add[3][3] , \PR_add[3][2] ,
         \PR_add[3][1] , \PR_add[3][0] , \PR_add[2][19] , \PR_add[2][18] ,
         \PR_add[2][17] , \PR_add[2][16] , \PR_add[2][15] , \PR_add[2][14] ,
         \PR_add[2][13] , \PR_add[2][12] , \PR_add[2][11] , \PR_add[2][10] ,
         \PR_add[2][9] , \PR_add[2][8] , \PR_add[2][7] , \PR_add[2][6] ,
         \PR_add[2][5] , \PR_add[2][4] , \PR_add[2][3] , \PR_add[2][2] ,
         \PR_add[1][19] , \PR_add[1][18] , \PR_add[1][17] , \PR_add[1][16] ,
         \PR_add[1][15] , \PR_add[1][14] , \PR_add[1][13] , \PR_add[1][12] ,
         \PR_add[1][11] , \PR_add[1][10] , \PR_add[1][9] , \PR_add[1][8] ,
         \PR_add[1][7] , \PR_add[1][6] , \PR_add[1][5] , \PR_add[1][4] ,
         \PR_add[1][3] , \PR_add[1][2] , \PR_add[1][1] , \PR_add[0][11] ,
         \PR_add[0][10] , \PR_add[0][9] , \PR_add[0][8] , \PR_add[0][7] ,
         \PR_add[0][6] , \PR_add[0][5] , \PR_add[0][4] , \PR_add[0][3] ,
         \PR_add[0][2] , \PR_add[0][1] , \PR_add[0][0] , N128, N129, N130,
         N131, N132, N133, N134, N135, N136, N137, N138, N139, N140, N148,
         N149, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159,
         N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170,
         N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181,
         N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192,
         N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203,
         N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214,
         N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225,
         N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236,
         N237, N238, N239, N240, N241, N242, N243, N244, N245, N246, N247,
         N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, N258,
         N259, N260, N261, N262, N263, N264, N265, N266, N267, N268, N269,
         N270, N271, N272, N273, N274, N275, N276, N277, N278, N279, N280,
         N281, N282, N283, N284, N285, N286, N287, N288, N289, N290, N291,
         N292, N293, N294, N295, N296, N297, N298, N299, N300, N301, N302,
         N303, N304, N305, N306, N307, N308, N309, N310, N311, N312, N313,
         N314, N315, N316, N317, N318, N319, N320, N321, N322, N323, N324,
         N325, N326, N327, N328, N329, N330, N331, N332, N333, N334, N335,
         N336, N337, N338, N339, N340, N341, N342, N343, N344, N345, N346,
         N347, N348, N349, N350, N351, N352, N353, N354, N355, N356, N357,
         N358, N359, N360, N361, N362, N363, N364, N365, N366, N367, N368,
         N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N401,
         N402, N403, N404, N405, N406, N407, N408, N409, N410, N411, N412,
         N413, N414, N415, N416, N417, N418, N419, N428, N429, N430, N431,
         N432, N433, N434, N435, N436, N437, N438, N439, N440, N448, N449,
         N450, N451, N452, N453, N454, N455, N456, N457, N458, N459, N460,
         N461, N462, N463, N464, N465, N466, N467, N468, N469, N470, N471,
         N472, N473, N474, N475, N476, N477, N478, N479, N480, N481, N482,
         N483, N484, N485, N486, N487, N488, N489, N490, N491, N492, N493,
         N494, N495, N496, N497, N498, N499, N500, N501, N502, N503, N504,
         N505, N506, N507, N508, N509, N510, N511, N512, N513, N514, N515,
         N516, N517, N518, N519, N520, N521, N522, N523, N524, N525, N526,
         N527, N528, N529, N530, N531, N532, N533, N534, N535, N536, N537,
         N538, N539, N540, N541, N542, N543, N544, N545, N546, N547, N548,
         N549, N550, N551, N552, N553, N554, N555, N556, N557, N558, N559,
         N560, N561, N562, N563, N564, N565, N566, N567, N568, N569, N570,
         N571, N572, N573, N574, N575, N576, N577, N578, N579, N580, N581,
         N582, N583, N584, N585, N586, N587, N588, N589, N590, N591, N592,
         N593, N594, N595, N596, N597, N598, N599, N600, N601, N602, N603,
         N604, N605, N606, N607, N608, N609, N610, N611, N612, N613, N614,
         N615, N616, N617, N618, N619, N620, N621, N622, N623, N624, N625,
         N626, N627, N628, N629, N630, N631, N632, N633, N634, N635, N636,
         N637, N638, N639, N640, N641, N642, N643, N644, N645, N646, N647,
         N648, N649, N650, N651, N652, N653, N654, N655, N656, N657, N658,
         N659, N660, N661, N662, N663, N664, N665, N666, N667, N668, N669,
         N670, N671, N672, N673, N674, N675, N676, N677, N678, N679, N680,
         N681, N682, N683, N684, N685, N686, N687, N688, N689, N690, N691,
         N692, N693, N694, N695, N704, N705, N706, N707, N708, N709, N710,
         N711, N712, N713, N714, N715, N716, N717, N718, N719, N728, N729,
         N730, N731, N732, N733, N734, N735, N744, N745, N746, N747, N748,
         N749, N750, N751, N752, N753, N754, N755, N756, N757, N758, N759,
         N768, N769, N770, N771, N772, N773, N774, N775, N784, N785, N786,
         N787, N788, N789, N790, N791, N792, N793, N794, N795, N796, N797,
         N798, N799, N800, N801, N802, N803, N804, N805, N806, N807, N808,
         N809, N810, N811, N812, N813, N814, N815, N816, N817, N818, N819,
         N820, N821, N822, N823, N824, N825, N826, N827, N828, N829, N830,
         N833, N834, N835, N836, N837, N838, N839, N840, N841, N842, N843,
         N844, N845, N846, N847, N848, N849, N850, N851, N852, N853, N854,
         N855, N856, N857, N858, N859, N860, N861, N862, N863, N864, N865,
         N866, N867, N868, N869, N870, N871, N872, N873, N874, N875, N876,
         N877, N878, N879, N880, N881, N884, N885, N886, N887, N888, N889,
         N890, N891, N892, N893, N894, N895, N896, N897, N898, N899, N900,
         N901, N902, N903, N904, N905, N906, N907, N908, N909, N910, N911,
         N912, N913, N914, N915, N916, N917, N918, N919, N920, N921, N922,
         N923, N924, N925, N926, N927, N928, N929, N930, N931, N932, N935,
         N936, N937, N938, N939, N940, N941, N942, N943, N944, N945, N946,
         N947, N948, N949, N950, N951, N952, N953, N954, N955, N956, N957,
         N958, N959, N960, N961, N962, N963, N964, N965, N966, N967, N968,
         N969, N970, N971, N972, m631, m633, m634, m635, m636, m637, m638,
         m639, m640, m641, m642, m643, m644, m645, m646, m647, m648, m649,
         m650, m651, m652, m653, m654, m655, m656, m657, m658, m659, m660,
         m661, m662, m663, m664, m665, m666, m667, m668, m669, m670, m673,
         m674, m675, m676, m677, m678, m679, m680, m681, m682, m683, m684,
         m685, m686, m687, m688, m689, m690, m691, m692, m693, m694, m695,
         m696, m697, m698, m699, m700, m701, m702, m703, m704, m705, m708,
         m709, m710, m711, m712, m713, m714, m715, m716, m717, m718, m719,
         m720, m721, m722, m723, m724, m725, m726, m727, m728, m729, m730,
         m731, m732, m733, m734, m735, m736, m737, m738, m739, m740, m743,
         m744, m745, m746, m747, m748, m749, m750, m751, m752, m753, m754,
         m755, m756, m757, m758, m759, m760, m761, m762, m763, m764, m765,
         m766, m767, m768, m769, m770, m771, m772, m773, m774, m775, m776,
         m777, m778, m779, m780, m781, m782, m784, m785, m786, m787, m788,
         m789, m790, m791, m792, m793, m794, m795, m796, m797, m798, m799,
         m800, m801, m802, m803, m804, m805, m806, m807, m808, m809, m810,
         m811, m812, m813, m814, m815, m816, m817, m818, m819, m820, m821,
         m822, m823, m824, m825, m826, m827, m828, m829, m830, m831, m832,
         m833, m834, m835, m836, m837, m838, m839, m840, m841, m842, m843,
         m844, m845, m846, m847, m848, m849, m850, m851, m852, m853, m854,
         m855, m856, m857, m858, m859, m860, m861, m862, m863, m864, m865,
         m866, m867, m868, m869, m870, m871, m872, m873, m874, m875, m876,
         m877, m878, m879, m880, m881, m882, m883, m884, m885, m886, m887,
         m888, m889, m890, m891, m892, m893, m894, m895, m896, m897, m898,
         m899, m900, m901, m902, m903, m904, m905, m906, m907, m908, m909,
         m910, m911, m912, m913, m914, m915, m916, m917, m918, m919, m920,
         m921, m922, m923, m924, m925, m926, m927, m928, m929, m930, m931,
         m932, m933, m934, m935, m936, m937, m938, m939, m940, m941, m942,
         m943, m944, m945, m946, m947, m948, m949, m950, m951, m952, m953,
         m954, m955, m956, m957, m958, m959, m960, m961, m962, m963, m964,
         m965, m966, m967, m968, m969, m970, m971, m972, m973, m974, m975,
         m976, m977, m978, m979, m980, m981, m982, m983, m984, m985, m986,
         m987, m988, m989, m990, m991, m992, m993, m994, m995, m996, m997,
         m998, m999, m1000, m1001, m1002, m1003, m1004, m1005, m1006, m1007,
         m1008, m1009, m1010, m1011, m1012, m1013, m1014, m1015, m1016, m1017,
         m1018, m1019, m1020, m1021, m1022, m1023, m1024, m1025, m1026, m1027,
         m1028, m1029, m1030, m1031, m1032, m1033, m1034, m1035, m1036, m1037,
         m1038, m1039, m1040, m1041, m1042, m1043, m1044, m1045, m1046, m1047,
         m1048, m1049, m1050, m1051, m1052, m1053, m1054, m1055, m1056, m1057,
         m1058, m1059, m1060, m1061, m1062, m1063, m1064, m1065, m1066, m1067,
         m1068, m1069, m1070, m1071, m1072, m1073, m1074, m1075, m1076, m1077,
         m1078, m1079, m1080, m1081, m1082, m1083, m1084, m1085, m1086, m1087,
         m1088, m1089, m1090, m1091, m1092, m1093, m1094, m1095, m1096, m1097,
         m1098, m1099, m1100, m1101, m1102, m1103, m1104, m1105, m1106, m1107,
         m1108, m1109, m1110, m1111, m1112, m1113, m1114, m1115, m1116, m1117,
         m1118, m1126, m1127, m1128, m1129, m1130, m1131, m1132, m1133, m1134,
         m1135, m1136, m1137, m1138, m1147, m1148, m1149, m1150, m1151, m1152,
         m1153, m1154, m1155, m1156, m1157, m1158, m1159, m1160, m1161, m1162,
         m1163, m1164, m1165, m1166, m1167, m1168, m1169, m1170, m1171, m1172,
         m1173, m1174, m1175, m1176, m1177, m1178, \mult_83/FS_1/P[0][0][1] ,
         \mult_83/FS_1/P[0][0][2] , \mult_83/FS_1/P[0][0][3] ,
         \mult_83/FS_1/P[0][1][1] , \mult_83/FS_1/P[0][1][2] ,
         \mult_83/FS_1/P[0][1][3] , \mult_83/FS_1/P[0][2][1] ,
         \mult_83/FS_1/TEMP_P[0][0][0] , \mult_83/FS_1/TEMP_P[0][1][0] ,
         \mult_83/FS_1/TEMP_P[0][2][0] , \mult_83/A2[9] , \mult_83/A1[0] ,
         \mult_83/A1[1] , \mult_83/A1[2] , \mult_83/A1[3] , \mult_83/A1[4] ,
         \mult_83/A1[5] , \mult_83/A1[6] , \mult_83/A1[7] , \mult_83/A1[8] ,
         \mult_83/ab[0][3] , \mult_83/ab[1][2] , \mult_83/ab[1][3] ,
         \mult_83/ab[2][2] , \mult_83/ab[2][3] , \mult_83/ab[3][2] ,
         \mult_83/ab[3][3] , \mult_83/ab[4][2] , \mult_83/ab[4][3] ,
         \mult_83/ab[5][2] , \mult_83/ab[5][3] , \mult_83/ab[6][2] ,
         \mult_83/ab[6][3] , \mult_83/ab[7][2] , \mult_83/ab[7][3] ,
         \mult_83/A_not[7] , \mult_80/FS_1/C[1][2][0] ,
         \mult_80/FS_1/P[0][0][1] , \mult_80/FS_1/P[0][0][2] ,
         \mult_80/FS_1/P[0][0][3] , \mult_80/FS_1/P[0][1][1] ,
         \mult_80/FS_1/P[0][1][2] , \mult_80/FS_1/P[0][1][3] ,
         \mult_80/FS_1/TEMP_P[0][0][0] , \mult_80/FS_1/TEMP_P[0][1][0] ,
         \mult_80/FS_1/TEMP_P[0][2][0] , \mult_80/FS_1/G[0][1][3] ,
         \mult_80/FS_1/G[1][0][1] , \mult_80/FS_1/G_n_int[0][1][3] ,
         \mult_80/FS_1/PG_int[0][2][0] , \mult_80/A2[7] , \mult_80/A2[8] ,
         \mult_80/A1[0] , \mult_80/A1[1] , \mult_80/A1[2] , \mult_80/A1[3] ,
         \mult_80/A1[4] , \mult_80/A1[5] , \mult_80/A1[6] , \mult_80/A1[7] ,
         \mult_80/ab[0][1] , \mult_80/ab[0][2] , \mult_80/ab[1][0] ,
         \mult_80/ab[1][1] , \mult_80/ab[1][2] , \mult_80/ab[2][0] ,
         \mult_80/ab[2][1] , \mult_80/ab[2][2] , \mult_80/ab[3][0] ,
         \mult_80/ab[3][1] , \mult_80/ab[3][2] , \mult_80/ab[4][0] ,
         \mult_80/ab[4][1] , \mult_80/ab[4][2] , \mult_80/ab[5][0] ,
         \mult_80/ab[5][1] , \mult_80/ab[5][2] , \mult_80/ab[6][0] ,
         \mult_80/ab[6][1] , \mult_80/ab[6][2] , \mult_80/ab[7][0] ,
         \mult_80/ab[7][1] , \mult_80/ab[7][2] , \mult_80/A_not[7] ,
         \mult_77/FS_1/P[0][0][1] , \mult_77/FS_1/P[0][0][2] ,
         \mult_77/FS_1/P[0][0][3] , \mult_77/FS_1/P[0][1][1] ,
         \mult_77/FS_1/P[0][1][2] , \mult_77/FS_1/P[0][1][3] ,
         \mult_77/FS_1/P[0][2][1] , \mult_77/FS_1/TEMP_P[0][0][0] ,
         \mult_77/FS_1/TEMP_P[0][1][0] , \mult_77/FS_1/TEMP_P[0][2][0] ,
         \mult_77/A2[9] , \mult_77/A1[0] , \mult_77/A1[1] , \mult_77/A1[2] ,
         \mult_77/A1[3] , \mult_77/A1[4] , \mult_77/A1[5] , \mult_77/A1[6] ,
         \mult_77/A1[7] , \mult_77/A1[8] , \mult_77/ab[0][3] ,
         \mult_77/ab[1][2] , \mult_77/ab[1][3] , \mult_77/ab[2][2] ,
         \mult_77/ab[2][3] , \mult_77/ab[3][2] , \mult_77/ab[3][3] ,
         \mult_77/ab[4][2] , \mult_77/ab[4][3] , \mult_77/ab[5][2] ,
         \mult_77/ab[5][3] , \mult_77/ab[6][2] , \mult_77/ab[6][3] ,
         \mult_77/ab[7][2] , \mult_77/ab[7][3] , \mult_77/A_not[7] ,
         \mult_76/FS_1/C[1][2][0] , \mult_76/FS_1/P[0][0][1] ,
         \mult_76/FS_1/P[0][0][2] , \mult_76/FS_1/P[0][0][3] ,
         \mult_76/FS_1/P[0][1][1] , \mult_76/FS_1/P[0][1][2] ,
         \mult_76/FS_1/P[0][1][3] , \mult_76/FS_1/TEMP_P[0][0][0] ,
         \mult_76/FS_1/TEMP_P[0][1][0] , \mult_76/FS_1/TEMP_P[0][2][0] ,
         \mult_76/FS_1/G[0][1][3] , \mult_76/FS_1/G[1][0][1] ,
         \mult_76/FS_1/G_n_int[0][1][3] , \mult_76/FS_1/PG_int[0][2][0] ,
         \mult_76/A2[7] , \mult_76/A1[0] , \mult_76/A1[1] , \mult_76/A1[2] ,
         \mult_76/A1[3] , \mult_76/A1[4] , \mult_76/A1[5] , \mult_76/A1[6] ,
         \mult_76/A1[7] , \mult_76/A1[8] , \mult_76/ab[0][3] ,
         \mult_76/ab[1][3] , \mult_76/ab[2][3] , \mult_76/ab[3][0] ,
         \mult_76/ab[3][3] , \mult_76/ab[4][0] , \mult_76/ab[4][3] ,
         \mult_76/ab[5][0] , \mult_76/ab[5][3] , \mult_76/ab[6][0] ,
         \mult_76/ab[7][0] , \mult_76/A_not[7] , \mult_74/FS_1/C[1][2][0] ,
         \mult_74/FS_1/P[0][0][1] , \mult_74/FS_1/P[0][0][2] ,
         \mult_74/FS_1/P[0][0][3] , \mult_74/FS_1/P[0][1][1] ,
         \mult_74/FS_1/P[0][1][2] , \mult_74/FS_1/P[0][1][3] ,
         \mult_74/FS_1/TEMP_P[0][0][0] , \mult_74/FS_1/TEMP_P[0][1][0] ,
         \mult_74/FS_1/TEMP_P[0][2][0] , \mult_74/FS_1/G[0][1][3] ,
         \mult_74/FS_1/G[1][0][1] , \mult_74/FS_1/G_n_int[0][1][3] ,
         \mult_74/FS_1/PG_int[0][2][0] , \mult_74/A2[7] , \mult_74/A2[8] ,
         \mult_74/A1[0] , \mult_74/A1[1] , \mult_74/A1[2] , \mult_74/A1[3] ,
         \mult_74/A1[4] , \mult_74/A1[5] , \mult_74/A1[6] , \mult_74/A1[7] ,
         \mult_74/ab[0][1] , \mult_74/ab[0][2] , \mult_74/ab[1][0] ,
         \mult_74/ab[1][1] , \mult_74/ab[1][2] , \mult_74/ab[2][0] ,
         \mult_74/ab[2][1] , \mult_74/ab[2][2] , \mult_74/ab[3][0] ,
         \mult_74/ab[3][1] , \mult_74/ab[3][2] , \mult_74/ab[4][0] ,
         \mult_74/ab[4][1] , \mult_74/ab[4][2] , \mult_74/ab[5][0] ,
         \mult_74/ab[5][1] , \mult_74/ab[5][2] , \mult_74/ab[6][0] ,
         \mult_74/ab[6][1] , \mult_74/ab[6][2] , \mult_74/ab[7][0] ,
         \mult_74/ab[7][1] , \mult_74/ab[7][2] , \mult_74/A_not[7] ,
         \mult_72/FS_1/P[0][0][1] , \mult_72/FS_1/P[0][0][2] ,
         \mult_72/FS_1/P[0][0][3] , \mult_72/FS_1/P[0][1][1] ,
         \mult_72/FS_1/P[0][1][2] , \mult_72/FS_1/P[0][1][3] ,
         \mult_72/FS_1/P[0][2][1] , \mult_72/FS_1/TEMP_P[0][0][0] ,
         \mult_72/FS_1/TEMP_P[0][1][0] , \mult_72/FS_1/TEMP_P[0][2][0] ,
         \mult_72/A2[9] , \mult_72/A1[0] , \mult_72/A1[1] , \mult_72/A1[2] ,
         \mult_72/A1[3] , \mult_72/A1[4] , \mult_72/A1[5] , \mult_72/A1[6] ,
         \mult_72/A1[7] , \mult_72/A1[8] , \mult_72/ab[0][3] ,
         \mult_72/ab[1][2] , \mult_72/ab[1][3] , \mult_72/ab[2][2] ,
         \mult_72/ab[2][3] , \mult_72/ab[3][2] , \mult_72/ab[3][3] ,
         \mult_72/ab[4][2] , \mult_72/ab[4][3] , \mult_72/ab[5][2] ,
         \mult_72/ab[5][3] , \mult_72/ab[6][2] , \mult_72/ab[6][3] ,
         \mult_72/ab[7][2] , \mult_72/ab[7][3] , \mult_72/A_not[7] ,
         \mult_71/FS_1/C[1][2][0] , \mult_71/FS_1/P[0][0][1] ,
         \mult_71/FS_1/P[0][0][2] , \mult_71/FS_1/P[0][0][3] ,
         \mult_71/FS_1/P[0][1][1] , \mult_71/FS_1/P[0][1][2] ,
         \mult_71/FS_1/P[0][1][3] , \mult_71/FS_1/TEMP_P[0][0][0] ,
         \mult_71/FS_1/TEMP_P[0][1][0] , \mult_71/FS_1/TEMP_P[0][2][0] ,
         \mult_71/FS_1/G[0][1][3] , \mult_71/FS_1/G[1][0][1] ,
         \mult_71/FS_1/G_n_int[0][1][3] , \mult_71/FS_1/PG_int[0][2][0] ,
         \mult_71/A2[7] , \mult_71/A1[0] , \mult_71/A1[1] , \mult_71/A1[2] ,
         \mult_71/A1[3] , \mult_71/A1[4] , \mult_71/A1[5] , \mult_71/A1[6] ,
         \mult_71/A1[7] , \mult_71/A1[8] , \mult_71/ab[0][3] ,
         \mult_71/ab[1][3] , \mult_71/ab[2][3] , \mult_71/ab[3][0] ,
         \mult_71/ab[3][3] , \mult_71/ab[4][0] , \mult_71/ab[4][3] ,
         \mult_71/ab[5][0] , \mult_71/ab[5][3] , \mult_71/ab[6][0] ,
         \mult_71/ab[7][0] , \mult_71/A_not[7] , \mult_69/FS_1/C[1][2][0] ,
         \mult_69/FS_1/P[0][0][1] , \mult_69/FS_1/P[0][0][2] ,
         \mult_69/FS_1/P[0][0][3] , \mult_69/FS_1/P[0][1][1] ,
         \mult_69/FS_1/P[0][1][2] , \mult_69/FS_1/P[0][1][3] ,
         \mult_69/FS_1/TEMP_P[0][0][0] , \mult_69/FS_1/TEMP_P[0][1][0] ,
         \mult_69/FS_1/TEMP_P[0][2][0] , \mult_69/FS_1/G[0][1][3] ,
         \mult_69/FS_1/G[1][0][1] , \mult_69/FS_1/G_n_int[0][1][3] ,
         \mult_69/FS_1/PG_int[0][2][0] , \mult_69/A2[7] , \mult_69/A2[8] ,
         \mult_69/A1[0] , \mult_69/A1[1] , \mult_69/A1[2] , \mult_69/A1[3] ,
         \mult_69/A1[4] , \mult_69/A1[5] , \mult_69/A1[6] , \mult_69/A1[7] ,
         \mult_69/ab[0][1] , \mult_69/ab[0][2] , \mult_69/ab[1][0] ,
         \mult_69/ab[1][1] , \mult_69/ab[1][2] , \mult_69/ab[2][0] ,
         \mult_69/ab[2][1] , \mult_69/ab[2][2] , \mult_69/ab[3][0] ,
         \mult_69/ab[3][1] , \mult_69/ab[3][2] , \mult_69/ab[4][0] ,
         \mult_69/ab[4][1] , \mult_69/ab[4][2] , \mult_69/ab[5][0] ,
         \mult_69/ab[5][1] , \mult_69/ab[5][2] , \mult_69/ab[6][0] ,
         \mult_69/ab[6][1] , \mult_69/ab[6][2] , \mult_69/ab[7][0] ,
         \mult_69/ab[7][1] , \mult_69/ab[7][2] , \mult_69/A_not[7] ,
         \mult_82/FS_1/C[1][2][0] , \mult_82/FS_1/P[0][0][1] ,
         \mult_82/FS_1/P[0][0][2] , \mult_82/FS_1/P[0][0][3] ,
         \mult_82/FS_1/P[0][1][1] , \mult_82/FS_1/P[0][1][2] ,
         \mult_82/FS_1/P[0][1][3] , \mult_82/FS_1/TEMP_P[0][0][0] ,
         \mult_82/FS_1/TEMP_P[0][1][0] , \mult_82/FS_1/TEMP_P[0][2][0] ,
         \mult_82/FS_1/G[0][1][3] , \mult_82/FS_1/G[1][0][1] ,
         \mult_82/FS_1/G_n_int[0][1][3] , \mult_82/FS_1/PG_int[0][2][0] ,
         \mult_82/A2[7] , \mult_82/A1[0] , \mult_82/A1[1] , \mult_82/A1[2] ,
         \mult_82/A1[3] , \mult_82/A1[4] , \mult_82/A1[5] , \mult_82/A1[6] ,
         \mult_82/A1[7] , \mult_82/A1[8] , \mult_82/ab[0][3] ,
         \mult_82/ab[1][3] , \mult_82/ab[2][3] , \mult_82/ab[3][0] ,
         \mult_82/ab[3][3] , \mult_82/ab[4][0] , \mult_82/ab[4][3] ,
         \mult_82/ab[5][0] , \mult_82/ab[5][3] , \mult_82/ab[6][0] ,
         \mult_82/ab[7][0] , \mult_82/A_not[7] , m1180, m1181, m1182, m1183,
         m1184, m1185, m1186, m1187, m1188, m1189, m1190, m1191, m1192, m1193,
         m1194, m1195, m1196, m1197, m1198, m1199, m1200, m1201, m1202, m1203,
         m1204, m1205, m1206, m1207, m1208, m1209, m1210, m1211, m1212, m1213,
         m1214, m1215, m1216, m1217, m1218, m1219, m1220, m1221, m1222, m1223,
         m1224, m1225, m1226, m1227, m1228, m1229, m1230, m1231, m1232, m1233,
         m1234, m1235, m1236, m1237, m1238, m1239, m1240, m1241, m1242, m1243,
         m1244, m1245, m1246, m1247, m1248, m1249, m1250, m1251, m1252, m1253,
         m1254, m1255, m1256, m1257, m1258, m1259, m1260, m1261, m1262, m1263,
         m1264, m1265, m1266, m1267, m1268, m1269, m1270, m1271, m1272, m1273,
         m1274, m1275, m1276, m1277, m1278, m1279, m1280, m1281, m1282, m1283,
         m1284, m1285, m1286, m1287, m1288, m1289, m1290, m1291, m1292, m1293,
         m1294, m1295, m1296, m1297, m1298, m1299, m1300, m1301, m1302, m1303,
         m1304, m1305, m1306, m1307, m1308, m1309, m1310, m1311, m1312, m1313,
         m1314, m1315, m1316, m1317, m1318, m1319, m1320, m1321, m1322, m1323,
         m1324, m1325, m1326, m1327, m1328, m1329, m1330, m1331, m1332, m1333,
         m1334, m1335, m1336, m1337, m1338, m1339, m1340, m1341, m1342, m1343,
         m1344, m1345, m1346, m1347, m1348, m1349, m1350, m1351, m1352, m1353,
         m1354, m1355, m1356, m1357, m1358, m1359, m1360, m1361, m1362, m1363,
         m1364, m1365, m1366, m1367, m1368, m1369, m1370, m1371, m1372, m1373,
         m1374, m1375, m1376, m1377, m1378, m1379, m1380, m1381, m1382, m1383,
         m1384, m1385, m1386, m1387, m1388, m1389, m1390, m1391, m1392, m1393,
         m1394, m1395, m1396, m1397, m1398, m1399, m1400, m1401, m1402, m1403,
         m1404, m1405, m1406, m1407, m1408, m1409, m1410, m1411, m1412, m1413,
         m1414, m1415, m1416, m1417, m1418, m1419, m1420, m1421, m1422, m1423,
         m1424, m1425, m1426, m1427, m1428, m1429, m1430, m1431, m1432, m1433,
         m1434, m1435, m1436, m1437, m1438, m1439, m1440, m1441, m1442, m1443,
         m1444, m1445, m1446, m1447, m1448, m1449, m1450, m1451, m1452, m1453,
         m1454, m1455, m1456, m1457, m1458, m1459, m1460, m1461, m1462, m1463,
         m1464, m1465, m1466, m1467, m1468, m1469, m1470, m1471, m1472, m1473,
         m1474, m1475, m1476, m1477, m1478, m1479, m1480, m1481, m1482, m1483,
         m1484, m1485, m1486, m1487, m1488, m1489, m1490, m1491, m1492, m1493,
         m1494, m1495, m1496, m1497, m1498, m1499, m1500, m1501, m1502, m1503,
         m1504, m1505, m1506, m1507, m1508, m1509, m1510, m1511, m1512, m1513,
         m1514, m1515, m1516, m1517, m1518, m1519, m1520, m1521, m1522, m1523,
         m1524, m1525, m1526, m1527, m1528, m1529, m1530, m1531, m1532, m1533,
         m1534, m1535, m1536, m1537, m1538, m1539, m1540, m1541, m1542, m1543,
         m1544, m1545, m1546, m1547, m1548, m1549, m1550, m1551, m1552, m1553,
         m1554, m1555, m1556, m1557, m1558, m1559, m1560, m1561, m1562, m1563,
         m1564, m1565, m1566, m1567, m1568, m1569, m1570, m1571, m1572, m1573,
         m1574, m1575, m1576, m1577, m1578, m1579, m1580, m1581, m1582, m1583,
         m1584, m1585, m1586, m1587, m1588, m1589, m1590, m1591, m1592, m1593,
         m1594, m1595, m1596, m1597, m1598, m1599, m1600, m1601, m1602, m1603,
         m1604, m1605, m1606, m1607, m1608, m1609, m1610, m1611, m1612, m1613,
         m1614, m1615, m1616, m1617, m1618, m1619, m1620, m1621, m1622, m1623,
         m1624, m1625, m1626, m1627, m1628, m1629, m1630, m1631, m1632, m1633,
         m1634, m1635, m1636, m1637, m1638, m1639, m1640, m1641, m1642, m1643,
         m1644, m1645, m1646, m1647, m1648, m1649, m1650, m1651, m1652, m1653,
         m1654, m1655, m1656, m1657, m1658, m1659, m1660, m1661, m1662, m1663,
         m1664, m1665, m1666, m1667, m1668, m1669, m1670, m1671, m1672, m1673,
         m1674, m1675, m1676, m1677, m1678, m1679, m1680, m1681, m1682, m1683,
         m1684, m1685, m1686, m1687, m1688, m1689, m1690, m1691, m1692, m1693,
         m1694, m1695, m1696, m1697, m1698, m1699, m1700, m1701, m1702, m1703,
         m1704, m1705, m1706, m1707, m1708, m1709, m1710, m1711, m1712, m1713,
         m1714, m1715, m1716, m1717, m1718, m1719, m1720, m1721, m1722, m1723,
         m1724, m1725, m1726, m1727, m1728, m1729, m1730, m1731, m1732, m1733,
         m1734, m1735, m1736, m1737, m1738, m1739, m1740, m1741, m1742, m1743,
         m1744, m1745, m1746, m1747, m1748, m1749, m1750, m1751, m1752, m1753,
         m1754, m1755, m1756, m1757, m1758, m1759, m1760, m1761, m1762, m1763,
         m1764, m1765, m1766, m1767, m1768, m1769, m1770, m1771, m1772, m1773,
         m1774, m1775, m1776, m1777, m1778, m1779, m1780, m1781, m1782, m1783,
         m1784, m1785, m1786, m1787, m1788, m1789, m1790, m1791, m1792, m1793,
         m1794, m1795, m1796, m1797, m1798, m1799, m1800, m1801, m1802, m1803,
         m1804, m1805, m1806, m1807, m1808, m1809, m1810, m1811, m1812, m1813,
         m1814, m1815, m1816, m1817, m1818, m1819, m1820, m1821, m1822, m1823,
         m1824, m1825, m1826, m1827, m1828, m1829, m1830, m1831, m1832, m1833,
         m1834, m1835, m1836, m1837, m1838, m1839, m1840, m1841, m1842, m1843,
         m1844, m1845, m1846, m1847, m1848, m1849, m1850, m1851, m1852, m1853,
         m1854, m1855, m1856, m1857, m1858, m1859, m1860, m1861, m1862, m1863,
         m1864, m1865, m1866, m1867, m1868, m1869, m1870, m1871, m1872, m1873,
         m1874, m1875, m1876, m1877, m1878, m1879, m1880, m1881, m1882, m1883,
         m1884, m1885, m1886, m1887, m1888, m1889, m1890, m1891, m1892, m1893,
         m1894, m1895, m1896, m1897, m1898, m1899, m1900, m1901, m1902, m1903,
         m1904, m1905, m1906, m1907, m1908, m1909, m1910, m1911, m1912, m1913,
         m1914, m1915, m1916, m1917, m1918, m1919, m1920, m1921, m1922, m1923,
         m1924, m1925, m1926, m1927, m1928, m1929, m1930, m1931, m1932, m1933,
         m1934, m1935, m1936, m1937, m1938, m1939, m1940, m1941, m1942, m1943,
         m1944, m1945, m1946, m1947, m1948, m1949, m1950, m1951, m1952, m1953,
         m1954, m1955, m1956, m1957, m1958, m1959, m1960, m1961, m1962, m1963,
         m1964, m1965, m1966, m1967, m1968, m1969, m1970, m1971, m1972, m1973,
         m1974, m1975, m1976, m1977, m1978, m1979, m1980, m1981, m1982, m1983,
         m1984, m1985, m1986, m1987, m1988, m1989, m1990, m1991, m1992, m1993,
         m1994, m1995, m1996, m1997, m1998, m1999, m2000, m2001, m2002, m2003,
         m2004, m2005, m2006, m2007, m2008, m2009, m2010, m2011, m2012, m2013,
         m2015, m2016, m2017, m2018, m2019, m2020, m2021, m2022, m2023, m2024,
         m2025, m2026, m2027, m2028, m2029, m2030, m2031, m2032, m2033, m2034,
         m2035, m2036, m2037, m2038, m2039, m2040, m2041, m2042, m2044, m2045,
         m2046, m2047, m2048, m2049, m2050, m2051, m2052, m2053, m2054, m2055,
         m2056, m2057, m2058, m2059, m2060, m2061, m2062, m2063, m2064, m2065,
         m2066, m2067, m2068, m2069, m2070, m2071, m2073, m2074, m2075, m2076,
         m2077, m2078, m2079, m2080, m2081, m2082, m2083, m2084, m2085, m2086,
         m2087, m2088, m2089, m2090, m2091, m2092, m2093, m2094, m2095, m2096,
         m2097, m2098, m2099, m2100, m2101, m2102, m2103, m2104, m2105, m2106,
         m2107, m2108, m2109, m2110, m2111, m2112, m2113, m2114, m2115, m2116,
         m2118, m2119, m2120, m2121, m2122, m2123, m2124, m2125, m2126, m2127,
         m2128, m2129, m2130, m2131, m2132, m2133, m2134, m2135, m2136, m2137,
         m2138, m2139, m2140, m2141, m2143, m2144, m2145, m2146, m2147, m2148,
         m2149, m2150, m2151, m2152, m2153, m2154, m2155, m2156, m2157, m2158,
         m2159, m2160, m2161, m2162, m2163, m2164, m2165, m2166, m2168, m2169,
         m2170, m2171, m2172, m2173, m2174, m2175, m2176, m2177, m2178, m2179,
         m2180, m2181, m2182, m2183, m2184, m2185, m2186, m2187, m2188, m2189,
         m2190, m2191, m2192, m2193, m2194, m2195, m2196, m2197, m2198, m2199,
         m2200, m2201, m2202, m2203, m2204, m2205, m2206, m2207, m2208, m2209,
         m2210, m2211, m2212, m2213, m2214, m2215, m2216, m2217, m2218, m2219,
         m2220, m2221, m2222, m2223, m2224, m2225, m2226, m2227, m2228, m2229,
         m2230, m2231, m2232, m2233, m2234, m2235, m2236, m2237, m2238, m2239,
         m2240, m2241, m2242, m2243, m2244, m2245, m2246, m2247, m2248, m2249,
         m2250, m2251, m2252, m2253, m2254, m2255, m2256, m2257, m2258, m2259,
         m2260, m2261, m2262, m2263, m2264, m2265, m2266, m2267, m2268, m2269,
         m2270, m2271, m2272, m2273, m2274, m2275, m2276, m2277, m2278, m2279,
         m2280, m2281, m2282, m2283, m2284, m2285, m2286, m2287, m2288, m2289,
         m2290, m2291, m2292, m2293, m2294, m2295, m2296, m2297, m2298, m2299,
         m2300, m2301, m2302, m2303, m2304, m2305, m2306, m2307, m2308, m2309,
         m2310, m2311, m2312, m2313, m2314, m2315, m2316, m2317, m2318, m2319,
         m2320, m2321, m2322, m2323, m2324, m2325, m2326, m2327, m2328, m2329,
         m2330, m2331, m2332, m2333, m2334, m2335, m2336, m2337, m2338, m2339,
         m2340, m2341, m2342, m2343, m2344, m2345, m2346, m2347, m2348, m2349,
         m2350, m2351, m2352, m2353, m2354, m2355, m2356, m2357, m2358, m2359,
         m2360, m2361, m2362, m2363, m2364, m2365, m2366, m2367, m2368, m2369,
         m2370, m2371, m2372, m2373, m2374, m2375, m2376, m2377, m2378, m2379,
         m2380, m2381, m2382, m2383, m2384, m2385, m2386, m2387, m2388, m2389,
         m2390, m2391, m2392, m2393, m2394, m2395, m2396, m2397, m2398, m2399,
         m2400, m2401, m2402, m2403, m2404, m2405, m2406, m2407, m2408, m2409,
         m2410, m2411, m2412, m2413, m2414, m2415, m2416, m2417, m2418, m2419,
         m2420, m2421, m2422, m2423, m2424, m2425, m2426, m2427, m2428, m2429,
         m2430, m2431, m2432, m2433, m2434, m2435, m2436, m2437, m2438, m2439,
         m2440, m2441, m2442, m2443, m2444, m2445, m2446, m2447, m2448, m2449,
         m2450, m2451, m2452, m2453, m2454, m2455, m2456, m2457, m2458, m2459,
         m2460, m2461, m2462, m2463, m2464, m2465, m2466, m2467, m2468, m2469,
         m2470, m2471, m2472, m2473, m2474, m2475, m2476, m2477, m2478, m2479,
         m2480, m2481, m2482, m2483, m2484, m2485, m2486, m2487, m2488, m2489,
         m2490, m2491, m2492, m2493, m2494, m2495, m2496, m2497, m2498, m2499,
         m2500, m2501, m2502, m2503, m2504, m2505, m2506, m2507, m2508, m2509,
         m2510, m2511, m2512, m2513, m2514, m2515, m2516, m2517, m2518, m2519,
         m2520, m2521, m2522, m2523, m2524, m2525, m2526, m2527, m2528, m2529,
         m2530, m2531, m2532, m2533, m2534, m2535, m2536, m2537, m2538, m2539,
         m2540, m2541, m2542, m2543, m2544, m2545, m2546, m2547, m2548, m2549,
         m2550, m2551, m2552, m2553, m2554, m2555, m2556, m2557, m2558, m2559,
         m2560, m2561, m2562, m2563, m2564, m2565, m2566, m2567, m2568, m2569,
         m2570, m2571, m2572, m2573, m2574, m2575, m2576, m2577, m2578, m2579,
         m2580, m2581, m2582, m2583, m2584, m2585, m2586, m2587, m2588, m2589,
         m2590, m2591, m2592, m2593, m2594, m2595, m2596, m2597, m2598, m2599,
         m2600;
  wire   [19:0] acc;
  wire   [6:0] \mult_83/A_notx ;
  wire   [6:0] \mult_80/A_notx ;
  wire   [6:0] \mult_77/A_notx ;
  wire   [6:0] \mult_76/A_notx ;
  wire   [6:0] \mult_74/A_notx ;
  wire   [6:0] \mult_72/A_notx ;
  wire   [6:0] \mult_71/A_notx ;
  wire   [6:0] \mult_69/A_notx ;
  wire   [6:0] \mult_82/A_notx ;

  Flip_Flop \PR_mul_reg[0][10]  ( .D(N810), .CLK(m1200), .R(1'b0), .Q(
        \PR_mul[0][10] ) );
  Flip_Flop \PR_mul_reg[0][9]  ( .D(N809), .CLK(m1201), .R(1'b0), .Q(
        \PR_mul[0][9] ) );
  Flip_Flop \PR_mul_reg[0][8]  ( .D(N808), .CLK(m1202), .R(1'b0), .Q(
        \PR_mul[0][8] ) );
  Flip_Flop \PR_mul_reg[0][7]  ( .D(N807), .CLK(m1204), .R(1'b0), .Q(
        \PR_mul[0][7] ) );
  Flip_Flop \PR_mul_reg[0][6]  ( .D(N806), .CLK(m1205), .R(1'b0), .Q(
        \PR_mul[0][6] ) );
  Flip_Flop \PR_mul_reg[0][5]  ( .D(N805), .CLK(m1207), .R(1'b0), .Q(
        \PR_mul[0][5] ) );
  Flip_Flop \PR_mul_reg[0][4]  ( .D(N804), .CLK(m1208), .R(1'b0), .Q(
        \PR_mul[0][4] ) );
  Flip_Flop \PR_mul_reg[0][3]  ( .D(N803), .CLK(m1210), .R(1'b0), .Q(
        \PR_mul[0][3] ) );
  Flip_Flop \PR_mul_reg[0][2]  ( .D(N802), .CLK(m1211), .R(1'b0), .Q(N110) );
  Flip_Flop \PR_mul_reg[0][1]  ( .D(N801), .CLK(m1212), .R(1'b0), .Q(N109) );
  Flip_Flop \PR_mul_reg[0][0]  ( .D(N800), .CLK(m1214), .R(1'b0), .Q(N108) );
  Flip_Flop \Samples_reg[0][7]  ( .D(N695), .CLK(m1218), .R(1'b0), .Q(
        \Samples[0][7] ) );
  Flip_Flop \PR_mul_reg[1][10]  ( .D(N818), .CLK(m1218), .R(1'b0), .Q(
        \PR_mul[1][10] ) );
  Flip_Flop \Samples_reg[1][7]  ( .D(N818), .CLK(m1218), .R(1'b0), .Q(
        \Samples[1][7] ) );
  Flip_Flop \Samples_reg[2][7]  ( .D(N711), .CLK(m1217), .R(1'b0), .Q(
        \Samples[2][7] ) );
  Flip_Flop \Samples_reg[3][7]  ( .D(N719), .CLK(m1217), .R(1'b0), .Q(
        \Samples[3][7] ) );
  Flip_Flop \PR_mul_reg[4][9]  ( .D(N850), .CLK(m1217), .R(1'b0), .Q(
        \PR_mul[4][9] ) );
  Flip_Flop \Samples_reg[4][7]  ( .D(N850), .CLK(m1217), .R(1'b0), .Q(
        \Samples[4][7] ) );
  Flip_Flop \Samples_reg[5][7]  ( .D(N735), .CLK(m1217), .R(1'b0), .Q(
        \Samples[5][7] ) );
  Flip_Flop \PR_mul_reg[6][10]  ( .D(N869), .CLK(m1216), .R(1'b0), .Q(
        \PR_mul[6][10] ) );
  Flip_Flop \Samples_reg[6][7]  ( .D(N869), .CLK(m1216), .R(1'b0), .Q(
        \Samples[6][7] ) );
  Flip_Flop \Samples_reg[7][7]  ( .D(N751), .CLK(m1216), .R(1'b0), .Q(
        \Samples[7][7] ) );
  Flip_Flop \Samples_reg[8][7]  ( .D(N759), .CLK(m1216), .R(1'b0), .Q(
        \Samples[8][7] ) );
  Flip_Flop \PR_mul_reg[9][9]  ( .D(N901), .CLK(m1215), .R(1'b0), .Q(
        \PR_mul[9][9] ) );
  Flip_Flop \Samples_reg[9][7]  ( .D(N901), .CLK(m1215), .R(1'b0), .Q(
        \Samples[9][7] ) );
  Flip_Flop \Samples_reg[10][7]  ( .D(N775), .CLK(m1215), .R(1'b0), .Q(
        \Samples[10][7] ) );
  Flip_Flop \PR_mul_reg[11][10]  ( .D(N920), .CLK(m1215), .R(1'b0), .Q(
        \PR_mul[11][10] ) );
  Flip_Flop \Samples_reg[11][7]  ( .D(N920), .CLK(m1215), .R(1'b0), .Q(
        \Samples[11][7] ) );
  Flip_Flop \Samples_reg[12][7]  ( .D(N791), .CLK(m1214), .R(1'b0), .Q(
        \Samples[12][7] ) );
  Flip_Flop \Samples_reg[13][7]  ( .D(N799), .CLK(m1214), .R(1'b0), .Q(
        \Samples[13][7] ) );
  Flip_Flop \PR_mul_reg[14][9]  ( .D(N952), .CLK(m1214), .R(1'b0), .Q(
        \PR_mul[14][9] ) );
  Flip_Flop \Samples_reg[0][6]  ( .D(N694), .CLK(m1220), .R(1'b0), .Q(
        \Samples[0][6] ) );
  Flip_Flop \PR_mul_reg[1][9]  ( .D(N817), .CLK(m1220), .R(1'b0), .Q(
        \PR_mul[1][9] ) );
  Flip_Flop \Samples_reg[1][6]  ( .D(N817), .CLK(m1220), .R(1'b0), .Q(
        \Samples[1][6] ) );
  Flip_Flop \Samples_reg[2][6]  ( .D(N710), .CLK(m1220), .R(1'b0), .Q(
        \Samples[2][6] ) );
  Flip_Flop \Samples_reg[3][6]  ( .D(N718), .CLK(m1220), .R(1'b0), .Q(
        \Samples[3][6] ) );
  Flip_Flop \PR_mul_reg[4][8]  ( .D(N849), .CLK(m1220), .R(1'b0), .Q(
        \PR_mul[4][8] ) );
  Flip_Flop \Samples_reg[4][6]  ( .D(N849), .CLK(m1220), .R(1'b0), .Q(
        \Samples[4][6] ) );
  Flip_Flop \Samples_reg[5][6]  ( .D(N734), .CLK(m1220), .R(1'b0), .Q(
        \Samples[5][6] ) );
  Flip_Flop \PR_mul_reg[6][9]  ( .D(N868), .CLK(m1220), .R(1'b0), .Q(
        \PR_mul[6][9] ) );
  Flip_Flop \Samples_reg[6][6]  ( .D(N868), .CLK(m1219), .R(1'b0), .Q(
        \Samples[6][6] ) );
  Flip_Flop \Samples_reg[7][6]  ( .D(N750), .CLK(m1219), .R(1'b0), .Q(
        \Samples[7][6] ) );
  Flip_Flop \Samples_reg[8][6]  ( .D(N758), .CLK(m1219), .R(1'b0), .Q(
        \Samples[8][6] ) );
  Flip_Flop \PR_mul_reg[9][8]  ( .D(N900), .CLK(m1219), .R(1'b0), .Q(
        \PR_mul[9][8] ) );
  Flip_Flop \Samples_reg[9][6]  ( .D(N900), .CLK(m1219), .R(1'b0), .Q(
        \Samples[9][6] ) );
  Flip_Flop \Samples_reg[10][6]  ( .D(N774), .CLK(m1219), .R(1'b0), .Q(
        \Samples[10][6] ) );
  Flip_Flop \PR_mul_reg[11][9]  ( .D(N919), .CLK(m1219), .R(1'b0), .Q(
        \PR_mul[11][9] ) );
  Flip_Flop \Samples_reg[11][6]  ( .D(N919), .CLK(m1219), .R(1'b0), .Q(
        \Samples[11][6] ) );
  Flip_Flop \Samples_reg[12][6]  ( .D(N790), .CLK(m1218), .R(1'b0), .Q(
        \Samples[12][6] ) );
  Flip_Flop \Samples_reg[13][6]  ( .D(N798), .CLK(m1218), .R(1'b0), .Q(
        \Samples[13][6] ) );
  Flip_Flop \PR_mul_reg[14][8]  ( .D(N951), .CLK(m1218), .R(1'b0), .Q(
        \PR_mul[14][8] ) );
  Flip_Flop \Samples_reg[0][5]  ( .D(N693), .CLK(m1223), .R(1'b0), .Q(
        \Samples[0][5] ) );
  Flip_Flop \PR_mul_reg[1][8]  ( .D(N816), .CLK(m1223), .R(1'b0), .Q(
        \PR_mul[1][8] ) );
  Flip_Flop \Samples_reg[1][5]  ( .D(N816), .CLK(m1223), .R(1'b0), .Q(
        \Samples[1][5] ) );
  Flip_Flop \Samples_reg[2][5]  ( .D(N709), .CLK(m1222), .R(1'b0), .Q(
        \Samples[2][5] ) );
  Flip_Flop \Samples_reg[3][5]  ( .D(N717), .CLK(m1222), .R(1'b0), .Q(
        \Samples[3][5] ) );
  Flip_Flop \PR_mul_reg[4][7]  ( .D(N848), .CLK(m1222), .R(1'b0), .Q(
        \PR_mul[4][7] ) );
  Flip_Flop \Samples_reg[4][5]  ( .D(N848), .CLK(m1222), .R(1'b0), .Q(
        \Samples[4][5] ) );
  Flip_Flop \Samples_reg[5][5]  ( .D(N733), .CLK(m1222), .R(1'b0), .Q(
        \Samples[5][5] ) );
  Flip_Flop \PR_mul_reg[6][8]  ( .D(N867), .CLK(m1222), .R(1'b0), .Q(
        \PR_mul[6][8] ) );
  Flip_Flop \Samples_reg[6][5]  ( .D(N867), .CLK(m1222), .R(1'b0), .Q(
        \Samples[6][5] ) );
  Flip_Flop \Samples_reg[7][5]  ( .D(N749), .CLK(m1222), .R(1'b0), .Q(
        \Samples[7][5] ) );
  Flip_Flop \Samples_reg[8][5]  ( .D(N757), .CLK(m1221), .R(1'b0), .Q(
        \Samples[8][5] ) );
  Flip_Flop \PR_mul_reg[9][7]  ( .D(N899), .CLK(m1221), .R(1'b0), .Q(
        \PR_mul[9][7] ) );
  Flip_Flop \Samples_reg[9][5]  ( .D(N899), .CLK(m1221), .R(1'b0), .Q(
        \Samples[9][5] ) );
  Flip_Flop \Samples_reg[10][5]  ( .D(N773), .CLK(m1221), .R(1'b0), .Q(
        \Samples[10][5] ) );
  Flip_Flop \PR_mul_reg[11][8]  ( .D(N918), .CLK(m1221), .R(1'b0), .Q(
        \PR_mul[11][8] ) );
  Flip_Flop \Samples_reg[11][5]  ( .D(N918), .CLK(m1221), .R(1'b0), .Q(
        \Samples[11][5] ) );
  Flip_Flop \Samples_reg[12][5]  ( .D(N789), .CLK(m1221), .R(1'b0), .Q(
        \Samples[12][5] ) );
  Flip_Flop \Samples_reg[13][5]  ( .D(N797), .CLK(m1221), .R(1'b0), .Q(
        \Samples[13][5] ) );
  Flip_Flop \PR_mul_reg[14][7]  ( .D(N950), .CLK(m1221), .R(1'b0), .Q(
        \PR_mul[14][7] ) );
  Flip_Flop \Samples_reg[0][4]  ( .D(N692), .CLK(m1225), .R(1'b0), .Q(
        \Samples[0][4] ) );
  Flip_Flop \PR_mul_reg[1][7]  ( .D(N815), .CLK(m1225), .R(1'b0), .Q(
        \PR_mul[1][7] ) );
  Flip_Flop \Samples_reg[1][4]  ( .D(N815), .CLK(m1225), .R(1'b0), .Q(
        \Samples[1][4] ) );
  Flip_Flop \Samples_reg[2][4]  ( .D(N708), .CLK(m1225), .R(1'b0), .Q(
        \Samples[2][4] ) );
  Flip_Flop \Samples_reg[3][4]  ( .D(N716), .CLK(m1225), .R(1'b0), .Q(
        \Samples[3][4] ) );
  Flip_Flop \PR_mul_reg[4][6]  ( .D(N847), .CLK(m1225), .R(1'b0), .Q(
        \PR_mul[4][6] ) );
  Flip_Flop \Samples_reg[4][4]  ( .D(N847), .CLK(m1224), .R(1'b0), .Q(
        \Samples[4][4] ) );
  Flip_Flop \Samples_reg[5][4]  ( .D(N732), .CLK(m1224), .R(1'b0), .Q(
        \Samples[5][4] ) );
  Flip_Flop \PR_mul_reg[6][7]  ( .D(N866), .CLK(m1224), .R(1'b0), .Q(
        \PR_mul[6][7] ) );
  Flip_Flop \Samples_reg[6][4]  ( .D(N866), .CLK(m1224), .R(1'b0), .Q(
        \Samples[6][4] ) );
  Flip_Flop \Samples_reg[7][4]  ( .D(N748), .CLK(m1224), .R(1'b0), .Q(
        \Samples[7][4] ) );
  Flip_Flop \Samples_reg[8][4]  ( .D(N756), .CLK(m1224), .R(1'b0), .Q(
        \Samples[8][4] ) );
  Flip_Flop \PR_mul_reg[9][6]  ( .D(N898), .CLK(m1224), .R(1'b0), .Q(
        \PR_mul[9][6] ) );
  Flip_Flop \Samples_reg[9][4]  ( .D(N898), .CLK(m1224), .R(1'b0), .Q(
        \Samples[9][4] ) );
  Flip_Flop \Samples_reg[10][4]  ( .D(N772), .CLK(m1223), .R(1'b0), .Q(
        \Samples[10][4] ) );
  Flip_Flop \PR_mul_reg[11][7]  ( .D(N917), .CLK(m1223), .R(1'b0), .Q(
        \PR_mul[11][7] ) );
  Flip_Flop \Samples_reg[11][4]  ( .D(N917), .CLK(m1223), .R(1'b0), .Q(
        \Samples[11][4] ) );
  Flip_Flop \Samples_reg[12][4]  ( .D(N788), .CLK(m1223), .R(1'b0), .Q(
        \Samples[12][4] ) );
  Flip_Flop \Samples_reg[13][4]  ( .D(N796), .CLK(m1223), .R(1'b0), .Q(
        \Samples[13][4] ) );
  Flip_Flop \PR_mul_reg[14][6]  ( .D(N949), .CLK(m1223), .R(1'b0), .Q(
        \PR_mul[14][6] ) );
  Flip_Flop \Samples_reg[0][3]  ( .D(N691), .CLK(m1227), .R(1'b0), .Q(
        \Samples[0][3] ) );
  Flip_Flop \PR_mul_reg[1][6]  ( .D(N814), .CLK(m1227), .R(1'b0), .Q(
        \PR_mul[1][6] ) );
  Flip_Flop \Samples_reg[1][3]  ( .D(N814), .CLK(m1227), .R(1'b0), .Q(
        \Samples[1][3] ) );
  Flip_Flop \Samples_reg[2][3]  ( .D(N707), .CLK(m1227), .R(1'b0), .Q(
        \Samples[2][3] ) );
  Flip_Flop \Samples_reg[3][3]  ( .D(N715), .CLK(m1227), .R(1'b0), .Q(
        \Samples[3][3] ) );
  Flip_Flop \PR_mul_reg[4][5]  ( .D(N846), .CLK(m1227), .R(1'b0), .Q(
        \PR_mul[4][5] ) );
  Flip_Flop \Samples_reg[4][3]  ( .D(N846), .CLK(m1227), .R(1'b0), .Q(
        \Samples[4][3] ) );
  Flip_Flop \Samples_reg[5][3]  ( .D(N731), .CLK(m1227), .R(1'b0), .Q(
        \Samples[5][3] ) );
  Flip_Flop \PR_mul_reg[6][6]  ( .D(N865), .CLK(m1227), .R(1'b0), .Q(
        \PR_mul[6][6] ) );
  Flip_Flop \Samples_reg[6][3]  ( .D(N865), .CLK(m1226), .R(1'b0), .Q(
        \Samples[6][3] ) );
  Flip_Flop \Samples_reg[7][3]  ( .D(N747), .CLK(m1226), .R(1'b0), .Q(
        \Samples[7][3] ) );
  Flip_Flop \Samples_reg[8][3]  ( .D(N755), .CLK(m1226), .R(1'b0), .Q(
        \Samples[8][3] ) );
  Flip_Flop \PR_mul_reg[9][5]  ( .D(N897), .CLK(m1226), .R(1'b0), .Q(
        \PR_mul[9][5] ) );
  Flip_Flop \Samples_reg[9][3]  ( .D(N897), .CLK(m1226), .R(1'b0), .Q(
        \Samples[9][3] ) );
  Flip_Flop \Samples_reg[10][3]  ( .D(N771), .CLK(m1226), .R(1'b0), .Q(
        \Samples[10][3] ) );
  Flip_Flop \PR_mul_reg[11][6]  ( .D(N916), .CLK(m1226), .R(1'b0), .Q(
        \PR_mul[11][6] ) );
  Flip_Flop \Samples_reg[11][3]  ( .D(N916), .CLK(m1226), .R(1'b0), .Q(
        \Samples[11][3] ) );
  Flip_Flop \Samples_reg[12][3]  ( .D(N787), .CLK(m1225), .R(1'b0), .Q(
        \Samples[12][3] ) );
  Flip_Flop \Samples_reg[13][3]  ( .D(N795), .CLK(m1225), .R(1'b0), .Q(
        \Samples[13][3] ) );
  Flip_Flop \PR_mul_reg[14][5]  ( .D(N948), .CLK(m1225), .R(1'b0), .Q(
        \PR_mul[14][5] ) );
  Flip_Flop \Samples_reg[0][2]  ( .D(N690), .CLK(m1230), .R(1'b0), .Q(
        \Samples[0][2] ) );
  Flip_Flop \PR_mul_reg[1][5]  ( .D(N813), .CLK(m1230), .R(1'b0), .Q(
        \PR_mul[1][5] ) );
  Flip_Flop \Samples_reg[1][2]  ( .D(N813), .CLK(m1230), .R(1'b0), .Q(
        \Samples[1][2] ) );
  Flip_Flop \Samples_reg[2][2]  ( .D(N706), .CLK(m1229), .R(1'b0), .Q(
        \Samples[2][2] ) );
  Flip_Flop \Samples_reg[3][2]  ( .D(N714), .CLK(m1229), .R(1'b0), .Q(
        \Samples[3][2] ) );
  Flip_Flop \PR_mul_reg[4][4]  ( .D(N845), .CLK(m1229), .R(1'b0), .Q(
        \PR_mul[4][4] ) );
  Flip_Flop \Samples_reg[4][2]  ( .D(N845), .CLK(m1229), .R(1'b0), .Q(
        \Samples[4][2] ) );
  Flip_Flop \Samples_reg[5][2]  ( .D(N730), .CLK(m1229), .R(1'b0), .Q(
        \Samples[5][2] ) );
  Flip_Flop \PR_mul_reg[6][5]  ( .D(N864), .CLK(m1229), .R(1'b0), .Q(
        \PR_mul[6][5] ) );
  Flip_Flop \Samples_reg[6][2]  ( .D(N864), .CLK(m1229), .R(1'b0), .Q(
        \Samples[6][2] ) );
  Flip_Flop \Samples_reg[7][2]  ( .D(N746), .CLK(m1229), .R(1'b0), .Q(
        \Samples[7][2] ) );
  Flip_Flop \Samples_reg[8][2]  ( .D(N754), .CLK(m1228), .R(1'b0), .Q(
        \Samples[8][2] ) );
  Flip_Flop \PR_mul_reg[9][4]  ( .D(N896), .CLK(m1228), .R(1'b0), .Q(
        \PR_mul[9][4] ) );
  Flip_Flop \Samples_reg[9][2]  ( .D(N896), .CLK(m1228), .R(1'b0), .Q(
        \Samples[9][2] ) );
  Flip_Flop \Samples_reg[10][2]  ( .D(N770), .CLK(m1228), .R(1'b0), .Q(
        \Samples[10][2] ) );
  Flip_Flop \PR_mul_reg[11][5]  ( .D(N915), .CLK(m1228), .R(1'b0), .Q(
        \PR_mul[11][5] ) );
  Flip_Flop \Samples_reg[11][2]  ( .D(N915), .CLK(m1228), .R(1'b0), .Q(
        \Samples[11][2] ) );
  Flip_Flop \Samples_reg[12][2]  ( .D(N786), .CLK(m1228), .R(1'b0), .Q(
        \Samples[12][2] ) );
  Flip_Flop \Samples_reg[13][2]  ( .D(N794), .CLK(m1228), .R(1'b0), .Q(
        \Samples[13][2] ) );
  Flip_Flop \PR_mul_reg[14][4]  ( .D(N947), .CLK(m1228), .R(1'b0), .Q(
        \PR_mul[14][4] ) );
  Flip_Flop \Samples_reg[0][1]  ( .D(N689), .CLK(m1232), .R(1'b0), .Q(
        \Samples[0][1] ) );
  Flip_Flop \PR_mul_reg[1][4]  ( .D(N812), .CLK(m1232), .R(1'b0), .Q(
        \PR_mul[1][4] ) );
  Flip_Flop \Samples_reg[1][1]  ( .D(N812), .CLK(m1232), .R(1'b0), .Q(
        \Samples[1][1] ) );
  Flip_Flop \Samples_reg[2][1]  ( .D(N705), .CLK(m1232), .R(1'b0), .Q(
        \Samples[2][1] ) );
  Flip_Flop \Samples_reg[3][1]  ( .D(N713), .CLK(m1232), .R(1'b0), .Q(
        \Samples[3][1] ) );
  Flip_Flop \PR_mul_reg[4][3]  ( .D(N844), .CLK(m1232), .R(1'b0), .Q(
        \PR_mul[4][3] ) );
  Flip_Flop \Samples_reg[4][1]  ( .D(N844), .CLK(m1231), .R(1'b0), .Q(
        \Samples[4][1] ) );
  Flip_Flop \Samples_reg[5][1]  ( .D(N729), .CLK(m1231), .R(1'b0), .Q(
        \Samples[5][1] ) );
  Flip_Flop \PR_mul_reg[6][4]  ( .D(N863), .CLK(m1231), .R(1'b0), .Q(
        \PR_mul[6][4] ) );
  Flip_Flop \Samples_reg[6][1]  ( .D(N863), .CLK(m1231), .R(1'b0), .Q(
        \Samples[6][1] ) );
  Flip_Flop \Samples_reg[7][1]  ( .D(N745), .CLK(m1231), .R(1'b0), .Q(
        \Samples[7][1] ) );
  Flip_Flop \Samples_reg[8][1]  ( .D(N753), .CLK(m1231), .R(1'b0), .Q(
        \Samples[8][1] ) );
  Flip_Flop \PR_mul_reg[9][3]  ( .D(N895), .CLK(m1231), .R(1'b0), .Q(
        \PR_mul[9][3] ) );
  Flip_Flop \Samples_reg[9][1]  ( .D(N895), .CLK(m1231), .R(1'b0), .Q(
        \Samples[9][1] ) );
  Flip_Flop \Samples_reg[10][1]  ( .D(N769), .CLK(m1230), .R(1'b0), .Q(
        \Samples[10][1] ) );
  Flip_Flop \PR_mul_reg[11][4]  ( .D(N914), .CLK(m1230), .R(1'b0), .Q(
        \PR_mul[11][4] ) );
  Flip_Flop \Samples_reg[11][1]  ( .D(N914), .CLK(m1230), .R(1'b0), .Q(
        \Samples[11][1] ) );
  Flip_Flop \Samples_reg[12][1]  ( .D(N785), .CLK(m1230), .R(1'b0), .Q(
        \Samples[12][1] ) );
  Flip_Flop \Samples_reg[13][1]  ( .D(N793), .CLK(m1230), .R(1'b0), .Q(
        \Samples[13][1] ) );
  Flip_Flop \PR_mul_reg[14][3]  ( .D(N946), .CLK(m1230), .R(1'b0), .Q(
        \PR_mul[14][3] ) );
  Flip_Flop \Samples_reg[0][0]  ( .D(N688), .CLK(m1234), .R(1'b0), .Q(
        \Samples[0][0] ) );
  Flip_Flop \PR_mul_reg[1][3]  ( .D(N811), .CLK(m1234), .R(1'b0), .Q(
        \PR_mul[1][3] ) );
  Flip_Flop \Samples_reg[1][0]  ( .D(N811), .CLK(m1234), .R(1'b0), .Q(
        \Samples[1][0] ) );
  Flip_Flop \PR_mul_reg[2][0]  ( .D(N819), .CLK(m1234), .R(1'b0), .Q(
        \PR_mul[2][0] ) );
  Flip_Flop \PR_mul_reg[2][1]  ( .D(N820), .CLK(m1232), .R(1'b0), .Q(
        \PR_mul[2][1] ) );
  Flip_Flop \PR_mul_reg[2][2]  ( .D(N821), .CLK(m1230), .R(1'b0), .Q(
        \PR_mul[2][2] ) );
  Flip_Flop \PR_mul_reg[2][3]  ( .D(N822), .CLK(m1227), .R(1'b0), .Q(
        \PR_mul[2][3] ) );
  Flip_Flop \PR_mul_reg[2][4]  ( .D(N823), .CLK(m1225), .R(1'b0), .Q(
        \PR_mul[2][4] ) );
  Flip_Flop \PR_mul_reg[2][5]  ( .D(N824), .CLK(m1223), .R(1'b0), .Q(
        \PR_mul[2][5] ) );
  Flip_Flop \PR_mul_reg[2][6]  ( .D(N825), .CLK(m1220), .R(1'b0), .Q(
        \PR_mul[2][6] ) );
  Flip_Flop \PR_mul_reg[2][7]  ( .D(N826), .CLK(m1218), .R(1'b0), .Q(
        \PR_mul[2][7] ) );
  Flip_Flop \PR_mul_reg[2][8]  ( .D(N827), .CLK(m1218), .R(1'b0), .Q(
        \PR_mul[2][8] ) );
  Flip_Flop \PR_mul_reg[2][9]  ( .D(N828), .CLK(m1218), .R(1'b0), .Q(
        \PR_mul[2][9] ) );
  Flip_Flop \PR_mul_reg[2][10]  ( .D(N829), .CLK(m1218), .R(1'b0), .Q(
        \PR_mul[2][10] ) );
  Flip_Flop \PR_mul_reg[2][11]  ( .D(N830), .CLK(m1218), .R(1'b0), .Q(
        \PR_mul[2][11] ) );
  Flip_Flop \Samples_reg[2][0]  ( .D(N704), .CLK(m1234), .R(1'b0), .Q(
        \Samples[2][0] ) );
  Flip_Flop \PR_mul_reg[3][2]  ( .D(N833), .CLK(m1234), .R(1'b0), .Q(
        \PR_mul[3][2] ) );
  Flip_Flop \PR_mul_reg[3][3]  ( .D(N834), .CLK(m1232), .R(1'b0), .Q(
        \PR_mul[3][3] ) );
  Flip_Flop \PR_mul_reg[3][4]  ( .D(N835), .CLK(m1229), .R(1'b0), .Q(
        \PR_mul[3][4] ) );
  Flip_Flop \PR_mul_reg[3][5]  ( .D(N836), .CLK(m1227), .R(1'b0), .Q(
        \PR_mul[3][5] ) );
  Flip_Flop \PR_mul_reg[3][6]  ( .D(N837), .CLK(m1225), .R(1'b0), .Q(
        \PR_mul[3][6] ) );
  Flip_Flop \PR_mul_reg[3][7]  ( .D(N838), .CLK(m1222), .R(1'b0), .Q(
        \PR_mul[3][7] ) );
  Flip_Flop \PR_mul_reg[3][8]  ( .D(N839), .CLK(m1220), .R(1'b0), .Q(
        \PR_mul[3][8] ) );
  Flip_Flop \PR_mul_reg[3][9]  ( .D(N840), .CLK(m1217), .R(1'b0), .Q(
        \PR_mul[3][9] ) );
  Flip_Flop \PR_mul_reg[3][10]  ( .D(N841), .CLK(m1217), .R(1'b0), .Q(
        \PR_mul[3][10] ) );
  Flip_Flop \PR_mul_reg[3][11]  ( .D(N842), .CLK(m1217), .R(1'b0), .Q(
        \PR_mul[3][11] ) );
  Flip_Flop \Samples_reg[3][0]  ( .D(N712), .CLK(m1234), .R(1'b0), .Q(
        \Samples[3][0] ) );
  Flip_Flop \PR_mul_reg[4][2]  ( .D(N843), .CLK(m1234), .R(1'b0), .Q(
        \PR_mul[4][2] ) );
  Flip_Flop \Samples_reg[4][0]  ( .D(N843), .CLK(m1234), .R(1'b0), .Q(
        \Samples[4][0] ) );
  Flip_Flop \PR_mul_reg[5][0]  ( .D(N851), .CLK(m1234), .R(1'b0), .Q(
        \PR_mul[5][0] ) );
  Flip_Flop \PR_mul_reg[5][1]  ( .D(N852), .CLK(m1231), .R(1'b0), .Q(
        \PR_mul[5][1] ) );
  Flip_Flop \PR_mul_reg[5][2]  ( .D(N853), .CLK(m1229), .R(1'b0), .Q(
        \PR_mul[5][2] ) );
  Flip_Flop \PR_mul_reg[5][3]  ( .D(N854), .CLK(m1227), .R(1'b0), .Q(
        \PR_mul[5][3] ) );
  Flip_Flop \PR_mul_reg[5][4]  ( .D(N855), .CLK(m1224), .R(1'b0), .Q(
        \PR_mul[5][4] ) );
  Flip_Flop \PR_mul_reg[5][5]  ( .D(N856), .CLK(m1222), .R(1'b0), .Q(
        \PR_mul[5][5] ) );
  Flip_Flop \PR_mul_reg[5][6]  ( .D(N857), .CLK(m1220), .R(1'b0), .Q(
        \PR_mul[5][6] ) );
  Flip_Flop \PR_mul_reg[5][7]  ( .D(N858), .CLK(m1217), .R(1'b0), .Q(
        \PR_mul[5][7] ) );
  Flip_Flop \PR_mul_reg[5][8]  ( .D(N859), .CLK(m1217), .R(1'b0), .Q(
        \PR_mul[5][8] ) );
  Flip_Flop \PR_mul_reg[5][9]  ( .D(N860), .CLK(m1217), .R(1'b0), .Q(
        \PR_mul[5][9] ) );
  Flip_Flop \PR_mul_reg[5][10]  ( .D(N861), .CLK(m1217), .R(1'b0), .Q(
        \PR_mul[5][10] ) );
  Flip_Flop \Samples_reg[5][0]  ( .D(N728), .CLK(m1234), .R(1'b0), .Q(
        \Samples[5][0] ) );
  Flip_Flop \PR_mul_reg[6][3]  ( .D(N862), .CLK(m1234), .R(1'b0), .Q(
        \PR_mul[6][3] ) );
  Flip_Flop \Samples_reg[6][0]  ( .D(N862), .CLK(m1233), .R(1'b0), .Q(
        \Samples[6][0] ) );
  Flip_Flop \PR_mul_reg[7][0]  ( .D(N870), .CLK(m1233), .R(1'b0), .Q(
        \PR_mul[7][0] ) );
  Flip_Flop \PR_mul_reg[7][1]  ( .D(N871), .CLK(m1231), .R(1'b0), .Q(
        \PR_mul[7][1] ) );
  Flip_Flop \PR_mul_reg[7][2]  ( .D(N872), .CLK(m1229), .R(1'b0), .Q(
        \PR_mul[7][2] ) );
  Flip_Flop \PR_mul_reg[7][3]  ( .D(N873), .CLK(m1226), .R(1'b0), .Q(
        \PR_mul[7][3] ) );
  Flip_Flop \PR_mul_reg[7][4]  ( .D(N874), .CLK(m1224), .R(1'b0), .Q(
        \PR_mul[7][4] ) );
  Flip_Flop \PR_mul_reg[7][5]  ( .D(N875), .CLK(m1222), .R(1'b0), .Q(
        \PR_mul[7][5] ) );
  Flip_Flop \PR_mul_reg[7][6]  ( .D(N876), .CLK(m1219), .R(1'b0), .Q(
        \PR_mul[7][6] ) );
  Flip_Flop \PR_mul_reg[7][7]  ( .D(N877), .CLK(m1216), .R(1'b0), .Q(
        \PR_mul[7][7] ) );
  Flip_Flop \PR_mul_reg[7][8]  ( .D(N878), .CLK(m1216), .R(1'b0), .Q(
        \PR_mul[7][8] ) );
  Flip_Flop \PR_mul_reg[7][9]  ( .D(N879), .CLK(m1216), .R(1'b0), .Q(
        \PR_mul[7][9] ) );
  Flip_Flop \PR_mul_reg[7][10]  ( .D(N880), .CLK(m1216), .R(1'b0), .Q(
        \PR_mul[7][10] ) );
  Flip_Flop \PR_mul_reg[7][11]  ( .D(N881), .CLK(m1216), .R(1'b0), .Q(
        \PR_mul[7][11] ) );
  Flip_Flop \Samples_reg[7][0]  ( .D(N744), .CLK(m1233), .R(1'b0), .Q(
        \Samples[7][0] ) );
  Flip_Flop \PR_mul_reg[8][2]  ( .D(N884), .CLK(m1233), .R(1'b0), .Q(
        \PR_mul[8][2] ) );
  Flip_Flop \PR_mul_reg[8][3]  ( .D(N885), .CLK(m1231), .R(1'b0), .Q(
        \PR_mul[8][3] ) );
  Flip_Flop \PR_mul_reg[8][4]  ( .D(N886), .CLK(m1229), .R(1'b0), .Q(
        \PR_mul[8][4] ) );
  Flip_Flop \PR_mul_reg[8][5]  ( .D(N887), .CLK(m1226), .R(1'b0), .Q(
        \PR_mul[8][5] ) );
  Flip_Flop \PR_mul_reg[8][6]  ( .D(N888), .CLK(m1224), .R(1'b0), .Q(
        \PR_mul[8][6] ) );
  Flip_Flop \PR_mul_reg[8][7]  ( .D(N889), .CLK(m1222), .R(1'b0), .Q(
        \PR_mul[8][7] ) );
  Flip_Flop \PR_mul_reg[8][8]  ( .D(N890), .CLK(m1219), .R(1'b0), .Q(
        \PR_mul[8][8] ) );
  Flip_Flop \PR_mul_reg[8][9]  ( .D(N891), .CLK(m1216), .R(1'b0), .Q(
        \PR_mul[8][9] ) );
  Flip_Flop \PR_mul_reg[8][10]  ( .D(N892), .CLK(m1216), .R(1'b0), .Q(
        \PR_mul[8][10] ) );
  Flip_Flop \PR_mul_reg[8][11]  ( .D(N893), .CLK(m1216), .R(1'b0), .Q(
        \PR_mul[8][11] ) );
  Flip_Flop \Samples_reg[8][0]  ( .D(N752), .CLK(m1233), .R(1'b0), .Q(
        \Samples[8][0] ) );
  Flip_Flop \PR_mul_reg[9][2]  ( .D(N894), .CLK(m1233), .R(1'b0), .Q(
        \PR_mul[9][2] ) );
  Flip_Flop \Samples_reg[9][0]  ( .D(N894), .CLK(m1233), .R(1'b0), .Q(
        \Samples[9][0] ) );
  Flip_Flop \PR_mul_reg[10][0]  ( .D(N902), .CLK(m1233), .R(1'b0), .Q(
        \PR_mul[10][0] ) );
  Flip_Flop \PR_mul_reg[10][1]  ( .D(N903), .CLK(m1231), .R(1'b0), .Q(
        \PR_mul[10][1] ) );
  Flip_Flop \PR_mul_reg[10][2]  ( .D(N904), .CLK(m1228), .R(1'b0), .Q(
        \PR_mul[10][2] ) );
  Flip_Flop \PR_mul_reg[10][3]  ( .D(N905), .CLK(m1226), .R(1'b0), .Q(
        \PR_mul[10][3] ) );
  Flip_Flop \PR_mul_reg[10][4]  ( .D(N906), .CLK(m1224), .R(1'b0), .Q(
        \PR_mul[10][4] ) );
  Flip_Flop \PR_mul_reg[10][5]  ( .D(N907), .CLK(m1221), .R(1'b0), .Q(
        \PR_mul[10][5] ) );
  Flip_Flop \PR_mul_reg[10][6]  ( .D(N908), .CLK(m1219), .R(1'b0), .Q(
        \PR_mul[10][6] ) );
  Flip_Flop \PR_mul_reg[10][7]  ( .D(N909), .CLK(m1215), .R(1'b0), .Q(
        \PR_mul[10][7] ) );
  Flip_Flop \PR_mul_reg[10][8]  ( .D(N910), .CLK(m1215), .R(1'b0), .Q(
        \PR_mul[10][8] ) );
  Flip_Flop \PR_mul_reg[10][9]  ( .D(N911), .CLK(m1215), .R(1'b0), .Q(
        \PR_mul[10][9] ) );
  Flip_Flop \PR_mul_reg[10][10]  ( .D(N912), .CLK(m1215), .R(1'b0), .Q(
        \PR_mul[10][10] ) );
  Flip_Flop \Samples_reg[10][0]  ( .D(N768), .CLK(m1233), .R(1'b0), .Q(
        \Samples[10][0] ) );
  Flip_Flop \PR_mul_reg[11][3]  ( .D(N913), .CLK(m1233), .R(1'b0), .Q(
        \PR_mul[11][3] ) );
  Flip_Flop \Samples_reg[11][0]  ( .D(N913), .CLK(m1233), .R(1'b0), .Q(
        \Samples[11][0] ) );
  Flip_Flop \PR_mul_reg[12][0]  ( .D(N921), .CLK(m1233), .R(1'b0), .Q(
        \PR_mul[12][0] ) );
  Flip_Flop \PR_mul_reg[12][1]  ( .D(N922), .CLK(m1230), .R(1'b0), .Q(
        \PR_mul[12][1] ) );
  Flip_Flop \PR_mul_reg[12][2]  ( .D(N923), .CLK(m1228), .R(1'b0), .Q(
        \PR_mul[12][2] ) );
  Flip_Flop \PR_mul_reg[12][3]  ( .D(N924), .CLK(m1226), .R(1'b0), .Q(
        \PR_mul[12][3] ) );
  Flip_Flop \PR_mul_reg[12][4]  ( .D(N925), .CLK(m1223), .R(1'b0), .Q(
        \PR_mul[12][4] ) );
  Flip_Flop \PR_mul_reg[12][5]  ( .D(N926), .CLK(m1221), .R(1'b0), .Q(
        \PR_mul[12][5] ) );
  Flip_Flop \PR_mul_reg[12][6]  ( .D(N927), .CLK(m1219), .R(1'b0), .Q(
        \PR_mul[12][6] ) );
  Flip_Flop \PR_mul_reg[12][7]  ( .D(N928), .CLK(m1215), .R(1'b0), .Q(
        \PR_mul[12][7] ) );
  Flip_Flop \PR_mul_reg[12][8]  ( .D(N929), .CLK(m1215), .R(1'b0), .Q(
        \PR_mul[12][8] ) );
  Flip_Flop \PR_mul_reg[12][9]  ( .D(N930), .CLK(m1214), .R(1'b0), .Q(
        \PR_mul[12][9] ) );
  Flip_Flop \PR_mul_reg[12][10]  ( .D(N931), .CLK(m1214), .R(1'b0), .Q(
        \PR_mul[12][10] ) );
  Flip_Flop \PR_mul_reg[12][11]  ( .D(N932), .CLK(m1215), .R(1'b0), .Q(
        \PR_mul[12][11] ) );
  Flip_Flop \Samples_reg[12][0]  ( .D(N784), .CLK(m1232), .R(1'b0), .Q(
        \Samples[12][0] ) );
  Flip_Flop \PR_mul_reg[13][2]  ( .D(N935), .CLK(m1232), .R(1'b0), .Q(
        \PR_mul[13][2] ) );
  Flip_Flop \PR_mul_reg[13][3]  ( .D(N936), .CLK(m1230), .R(1'b0), .Q(
        \PR_mul[13][3] ) );
  Flip_Flop \PR_mul_reg[13][4]  ( .D(N937), .CLK(m1228), .R(1'b0), .Q(
        \PR_mul[13][4] ) );
  Flip_Flop \PR_mul_reg[13][5]  ( .D(N938), .CLK(m1225), .R(1'b0), .Q(
        \PR_mul[13][5] ) );
  Flip_Flop \PR_mul_reg[13][6]  ( .D(N939), .CLK(m1223), .R(1'b0), .Q(
        \PR_mul[13][6] ) );
  Flip_Flop \PR_mul_reg[13][7]  ( .D(N940), .CLK(m1221), .R(1'b0), .Q(
        \PR_mul[13][7] ) );
  Flip_Flop \PR_mul_reg[13][8]  ( .D(N941), .CLK(m1218), .R(1'b0), .Q(
        \PR_mul[13][8] ) );
  Flip_Flop \PR_mul_reg[13][9]  ( .D(N942), .CLK(m1214), .R(1'b0), .Q(
        \PR_mul[13][9] ) );
  Flip_Flop \PR_mul_reg[13][10]  ( .D(N943), .CLK(m1214), .R(1'b0), .Q(
        \PR_mul[13][10] ) );
  Flip_Flop \PR_mul_reg[13][11]  ( .D(N944), .CLK(m1214), .R(1'b0), .Q(
        \PR_mul[13][11] ) );
  Flip_Flop \Samples_reg[13][0]  ( .D(N792), .CLK(m1232), .R(1'b0), .Q(
        \Samples[13][0] ) );
  Flip_Flop \PR_mul_reg[14][2]  ( .D(N945), .CLK(m1232), .R(1'b0), .Q(
        \PR_mul[14][2] ) );
  Flip_Flop \PR_add_reg[0][11]  ( .D(N419), .CLK(m1200), .R(1'b0), .Q(
        \PR_add[0][11] ) );
  Flip_Flop \PR_add_reg[0][10]  ( .D(N418), .CLK(m1199), .R(1'b0), .Q(
        \PR_add[0][10] ) );
  Flip_Flop \PR_add_reg[0][9]  ( .D(N417), .CLK(m1201), .R(1'b0), .Q(
        \PR_add[0][9] ) );
  Flip_Flop \PR_add_reg[0][8]  ( .D(N416), .CLK(m1202), .R(1'b0), .Q(
        \PR_add[0][8] ) );
  Flip_Flop \PR_add_reg[0][7]  ( .D(N415), .CLK(m1204), .R(1'b0), .Q(
        \PR_add[0][7] ) );
  Flip_Flop \PR_add_reg[0][6]  ( .D(N414), .CLK(m1205), .R(1'b0), .Q(
        \PR_add[0][6] ) );
  Flip_Flop \PR_add_reg[0][5]  ( .D(N413), .CLK(m1207), .R(1'b0), .Q(
        \PR_add[0][5] ) );
  Flip_Flop \PR_add_reg[0][4]  ( .D(N412), .CLK(m1208), .R(1'b0), .Q(
        \PR_add[0][4] ) );
  Flip_Flop \PR_add_reg[0][3]  ( .D(N411), .CLK(m1209), .R(1'b0), .Q(
        \PR_add[0][3] ) );
  Flip_Flop \PR_add_reg[0][2]  ( .D(N410), .CLK(m1211), .R(1'b0), .Q(
        \PR_add[0][2] ) );
  Flip_Flop \PR_add_reg[0][1]  ( .D(N409), .CLK(m1212), .R(1'b0), .Q(
        \PR_add[0][1] ) );
  Flip_Flop \PR_add_reg[0][0]  ( .D(N408), .CLK(m1214), .R(1'b0), .Q(
        \PR_add[0][0] ) );
  Flip_Flop \PR_add_reg[1][0]  ( .D(N428), .CLK(m1214), .R(1'b0), .Q(N148) );
  Flip_Flop \PR_add_reg[1][1]  ( .D(N429), .CLK(m1212), .R(1'b0), .Q(
        \PR_add[1][1] ) );
  Flip_Flop \PR_add_reg[1][2]  ( .D(N430), .CLK(m1211), .R(1'b0), .Q(
        \PR_add[1][2] ) );
  Flip_Flop \PR_add_reg[1][3]  ( .D(N431), .CLK(m1209), .R(1'b0), .Q(
        \PR_add[1][3] ) );
  Flip_Flop \PR_add_reg[1][4]  ( .D(N432), .CLK(m1208), .R(1'b0), .Q(
        \PR_add[1][4] ) );
  Flip_Flop \PR_add_reg[1][5]  ( .D(N433), .CLK(m1207), .R(1'b0), .Q(
        \PR_add[1][5] ) );
  Flip_Flop \PR_add_reg[1][6]  ( .D(N434), .CLK(m1205), .R(1'b0), .Q(
        \PR_add[1][6] ) );
  Flip_Flop \PR_add_reg[1][7]  ( .D(N435), .CLK(m1204), .R(1'b0), .Q(
        \PR_add[1][7] ) );
  Flip_Flop \PR_add_reg[1][8]  ( .D(N436), .CLK(m1202), .R(1'b0), .Q(
        \PR_add[1][8] ) );
  Flip_Flop \PR_add_reg[1][9]  ( .D(N437), .CLK(m1201), .R(1'b0), .Q(
        \PR_add[1][9] ) );
  Flip_Flop \PR_add_reg[1][10]  ( .D(N438), .CLK(m1199), .R(1'b0), .Q(
        \PR_add[1][10] ) );
  Flip_Flop \PR_add_reg[1][11]  ( .D(N439), .CLK(m1199), .R(1'b0), .Q(
        \PR_add[1][11] ) );
  Flip_Flop \PR_add_reg[1][12]  ( .D(N440), .CLK(m1199), .R(1'b0), .Q(
        \PR_add[1][12] ) );
  Flip_Flop \PR_add_reg[1][13]  ( .D(1'b0), .CLK(m1235), .R(1'b0), .Q(
        \PR_add[1][13] ) );
  Flip_Flop \PR_add_reg[1][14]  ( .D(1'b0), .CLK(m1235), .R(1'b0), .Q(
        \PR_add[1][14] ) );
  Flip_Flop \PR_add_reg[1][15]  ( .D(1'b0), .CLK(m1235), .R(1'b0), .Q(
        \PR_add[1][15] ) );
  Flip_Flop \PR_add_reg[1][16]  ( .D(1'b0), .CLK(m1235), .R(1'b0), .Q(
        \PR_add[1][16] ) );
  Flip_Flop \PR_add_reg[1][17]  ( .D(1'b0), .CLK(m1235), .R(1'b0), .Q(
        \PR_add[1][17] ) );
  Flip_Flop \PR_add_reg[1][18]  ( .D(1'b0), .CLK(m1235), .R(1'b0), .Q(
        \PR_add[1][18] ) );
  Flip_Flop \PR_add_reg[1][19]  ( .D(1'b0), .CLK(m1235), .R(1'b0), .Q(
        \PR_add[1][19] ) );
  Flip_Flop \PR_add_reg[2][0]  ( .D(N448), .CLK(m1214), .R(1'b0), .Q(N168) );
  Flip_Flop \PR_add_reg[2][1]  ( .D(N449), .CLK(m1212), .R(1'b0), .Q(N169) );
  Flip_Flop \PR_add_reg[2][2]  ( .D(N450), .CLK(m1211), .R(1'b0), .Q(
        \PR_add[2][2] ) );
  Flip_Flop \PR_add_reg[2][3]  ( .D(N451), .CLK(m1209), .R(1'b0), .Q(
        \PR_add[2][3] ) );
  Flip_Flop \PR_add_reg[2][4]  ( .D(N452), .CLK(m1208), .R(1'b0), .Q(
        \PR_add[2][4] ) );
  Flip_Flop \PR_add_reg[2][5]  ( .D(N453), .CLK(m1206), .R(1'b0), .Q(
        \PR_add[2][5] ) );
  Flip_Flop \PR_add_reg[2][6]  ( .D(N454), .CLK(m1205), .R(1'b0), .Q(
        \PR_add[2][6] ) );
  Flip_Flop \PR_add_reg[2][7]  ( .D(N455), .CLK(m1204), .R(1'b0), .Q(
        \PR_add[2][7] ) );
  Flip_Flop \PR_add_reg[2][8]  ( .D(N456), .CLK(m1202), .R(1'b0), .Q(
        \PR_add[2][8] ) );
  Flip_Flop \PR_add_reg[2][9]  ( .D(N457), .CLK(m1201), .R(1'b0), .Q(
        \PR_add[2][9] ) );
  Flip_Flop \PR_add_reg[2][10]  ( .D(N458), .CLK(m1198), .R(1'b0), .Q(
        \PR_add[2][10] ) );
  Flip_Flop \PR_add_reg[2][11]  ( .D(N459), .CLK(m1198), .R(1'b0), .Q(
        \PR_add[2][11] ) );
  Flip_Flop \PR_add_reg[2][12]  ( .D(N460), .CLK(m1199), .R(1'b0), .Q(
        \PR_add[2][12] ) );
  Flip_Flop \PR_add_reg[2][13]  ( .D(N461), .CLK(m1199), .R(1'b0), .Q(
        \PR_add[2][13] ) );
  Flip_Flop \PR_add_reg[2][14]  ( .D(N462), .CLK(m1199), .R(1'b0), .Q(
        \PR_add[2][14] ) );
  Flip_Flop \PR_add_reg[2][15]  ( .D(N463), .CLK(m1199), .R(1'b0), .Q(
        \PR_add[2][15] ) );
  Flip_Flop \PR_add_reg[2][16]  ( .D(N464), .CLK(m1199), .R(1'b0), .Q(
        \PR_add[2][16] ) );
  Flip_Flop \PR_add_reg[2][17]  ( .D(N465), .CLK(m1199), .R(1'b0), .Q(
        \PR_add[2][17] ) );
  Flip_Flop \PR_add_reg[2][18]  ( .D(N466), .CLK(m1199), .R(1'b0), .Q(
        \PR_add[2][18] ) );
  Flip_Flop \PR_add_reg[2][19]  ( .D(N467), .CLK(m1199), .R(1'b0), .Q(
        \PR_add[2][19] ) );
  Flip_Flop \PR_add_reg[3][0]  ( .D(N468), .CLK(m1213), .R(1'b0), .Q(
        \PR_add[3][0] ) );
  Flip_Flop \PR_add_reg[3][1]  ( .D(N469), .CLK(m1212), .R(1'b0), .Q(
        \PR_add[3][1] ) );
  Flip_Flop \PR_add_reg[3][2]  ( .D(N470), .CLK(m1211), .R(1'b0), .Q(
        \PR_add[3][2] ) );
  Flip_Flop \PR_add_reg[3][3]  ( .D(N471), .CLK(m1209), .R(1'b0), .Q(
        \PR_add[3][3] ) );
  Flip_Flop \PR_add_reg[3][4]  ( .D(N472), .CLK(m1208), .R(1'b0), .Q(
        \PR_add[3][4] ) );
  Flip_Flop \PR_add_reg[3][5]  ( .D(N473), .CLK(m1206), .R(1'b0), .Q(
        \PR_add[3][5] ) );
  Flip_Flop \PR_add_reg[3][6]  ( .D(N474), .CLK(m1205), .R(1'b0), .Q(
        \PR_add[3][6] ) );
  Flip_Flop \PR_add_reg[3][7]  ( .D(N475), .CLK(m1204), .R(1'b0), .Q(
        \PR_add[3][7] ) );
  Flip_Flop \PR_add_reg[3][8]  ( .D(N476), .CLK(m1202), .R(1'b0), .Q(
        \PR_add[3][8] ) );
  Flip_Flop \PR_add_reg[3][9]  ( .D(N477), .CLK(m1201), .R(1'b0), .Q(
        \PR_add[3][9] ) );
  Flip_Flop \PR_add_reg[3][10]  ( .D(N478), .CLK(m1198), .R(1'b0), .Q(
        \PR_add[3][10] ) );
  Flip_Flop \PR_add_reg[3][11]  ( .D(N479), .CLK(m1198), .R(1'b0), .Q(
        \PR_add[3][11] ) );
  Flip_Flop \PR_add_reg[3][12]  ( .D(N480), .CLK(m1196), .R(1'b0), .Q(
        \PR_add[3][12] ) );
  Flip_Flop \PR_add_reg[3][13]  ( .D(N481), .CLK(m1195), .R(1'b0), .Q(
        \PR_add[3][13] ) );
  Flip_Flop \PR_add_reg[3][14]  ( .D(N482), .CLK(m1195), .R(1'b0), .Q(
        \PR_add[3][14] ) );
  Flip_Flop \PR_add_reg[3][15]  ( .D(N483), .CLK(m1195), .R(1'b0), .Q(
        \PR_add[3][15] ) );
  Flip_Flop \PR_add_reg[3][16]  ( .D(N484), .CLK(m1195), .R(1'b0), .Q(
        \PR_add[3][16] ) );
  Flip_Flop \PR_add_reg[3][17]  ( .D(N485), .CLK(m1195), .R(1'b0), .Q(
        \PR_add[3][17] ) );
  Flip_Flop \PR_add_reg[3][18]  ( .D(N486), .CLK(m1195), .R(1'b0), .Q(
        \PR_add[3][18] ) );
  Flip_Flop \PR_add_reg[3][19]  ( .D(N487), .CLK(m1195), .R(1'b0), .Q(
        \PR_add[3][19] ) );
  Flip_Flop \PR_add_reg[4][0]  ( .D(N488), .CLK(m1213), .R(1'b0), .Q(N208) );
  Flip_Flop \PR_add_reg[4][1]  ( .D(N489), .CLK(m1212), .R(1'b0), .Q(N209) );
  Flip_Flop \PR_add_reg[4][2]  ( .D(N490), .CLK(m1211), .R(1'b0), .Q(N210) );
  Flip_Flop \PR_add_reg[4][3]  ( .D(N491), .CLK(m1209), .R(1'b0), .Q(
        \PR_add[4][3] ) );
  Flip_Flop \PR_add_reg[4][4]  ( .D(N492), .CLK(m1208), .R(1'b0), .Q(
        \PR_add[4][4] ) );
  Flip_Flop \PR_add_reg[4][5]  ( .D(N493), .CLK(m1206), .R(1'b0), .Q(
        \PR_add[4][5] ) );
  Flip_Flop \PR_add_reg[4][6]  ( .D(N494), .CLK(m1205), .R(1'b0), .Q(
        \PR_add[4][6] ) );
  Flip_Flop \PR_add_reg[4][7]  ( .D(N495), .CLK(m1203), .R(1'b0), .Q(
        \PR_add[4][7] ) );
  Flip_Flop \PR_add_reg[4][8]  ( .D(N496), .CLK(m1202), .R(1'b0), .Q(
        \PR_add[4][8] ) );
  Flip_Flop \PR_add_reg[4][9]  ( .D(N497), .CLK(m1201), .R(1'b0), .Q(
        \PR_add[4][9] ) );
  Flip_Flop \PR_add_reg[4][10]  ( .D(N498), .CLK(m1198), .R(1'b0), .Q(
        \PR_add[4][10] ) );
  Flip_Flop \PR_add_reg[4][11]  ( .D(N499), .CLK(m1198), .R(1'b0), .Q(
        \PR_add[4][11] ) );
  Flip_Flop \PR_add_reg[4][12]  ( .D(N500), .CLK(m1196), .R(1'b0), .Q(
        \PR_add[4][12] ) );
  Flip_Flop \PR_add_reg[4][13]  ( .D(N501), .CLK(m1194), .R(1'b0), .Q(
        \PR_add[4][13] ) );
  Flip_Flop \PR_add_reg[4][14]  ( .D(N502), .CLK(m1193), .R(1'b0), .Q(
        \PR_add[4][14] ) );
  Flip_Flop \PR_add_reg[4][15]  ( .D(N503), .CLK(m1193), .R(1'b0), .Q(
        \PR_add[4][15] ) );
  Flip_Flop \PR_add_reg[4][16]  ( .D(N504), .CLK(m1193), .R(1'b0), .Q(
        \PR_add[4][16] ) );
  Flip_Flop \PR_add_reg[4][17]  ( .D(N505), .CLK(m1193), .R(1'b0), .Q(
        \PR_add[4][17] ) );
  Flip_Flop \PR_add_reg[4][18]  ( .D(N506), .CLK(m1193), .R(1'b0), .Q(
        \PR_add[4][18] ) );
  Flip_Flop \PR_add_reg[4][19]  ( .D(N507), .CLK(m1193), .R(1'b0), .Q(
        \PR_add[4][19] ) );
  Flip_Flop \PR_add_reg[5][0]  ( .D(N508), .CLK(m1213), .R(1'b0), .Q(
        \PR_add[5][0] ) );
  Flip_Flop \PR_add_reg[5][1]  ( .D(N509), .CLK(m1212), .R(1'b0), .Q(
        \PR_add[5][1] ) );
  Flip_Flop \PR_add_reg[5][2]  ( .D(N510), .CLK(m1210), .R(1'b0), .Q(
        \PR_add[5][2] ) );
  Flip_Flop \PR_add_reg[5][3]  ( .D(N511), .CLK(m1209), .R(1'b0), .Q(
        \PR_add[5][3] ) );
  Flip_Flop \PR_add_reg[5][4]  ( .D(N512), .CLK(m1208), .R(1'b0), .Q(
        \PR_add[5][4] ) );
  Flip_Flop \PR_add_reg[5][5]  ( .D(N513), .CLK(m1206), .R(1'b0), .Q(
        \PR_add[5][5] ) );
  Flip_Flop \PR_add_reg[5][6]  ( .D(N514), .CLK(m1205), .R(1'b0), .Q(
        \PR_add[5][6] ) );
  Flip_Flop \PR_add_reg[5][7]  ( .D(N515), .CLK(m1203), .R(1'b0), .Q(
        \PR_add[5][7] ) );
  Flip_Flop \PR_add_reg[5][8]  ( .D(N516), .CLK(m1202), .R(1'b0), .Q(
        \PR_add[5][8] ) );
  Flip_Flop \PR_add_reg[5][9]  ( .D(N517), .CLK(m1201), .R(1'b0), .Q(
        \PR_add[5][9] ) );
  Flip_Flop \PR_add_reg[5][10]  ( .D(N518), .CLK(m1198), .R(1'b0), .Q(
        \PR_add[5][10] ) );
  Flip_Flop \PR_add_reg[5][11]  ( .D(N519), .CLK(m1198), .R(1'b0), .Q(
        \PR_add[5][11] ) );
  Flip_Flop \PR_add_reg[5][12]  ( .D(N520), .CLK(m1196), .R(1'b0), .Q(
        \PR_add[5][12] ) );
  Flip_Flop \PR_add_reg[5][13]  ( .D(N521), .CLK(m1194), .R(1'b0), .Q(
        \PR_add[5][13] ) );
  Flip_Flop \PR_add_reg[5][14]  ( .D(N522), .CLK(m1193), .R(1'b0), .Q(
        \PR_add[5][14] ) );
  Flip_Flop \PR_add_reg[5][15]  ( .D(N523), .CLK(m1192), .R(1'b0), .Q(
        \PR_add[5][15] ) );
  Flip_Flop \PR_add_reg[5][16]  ( .D(N524), .CLK(m1191), .R(1'b0), .Q(
        \PR_add[5][16] ) );
  Flip_Flop \PR_add_reg[5][17]  ( .D(N525), .CLK(m1191), .R(1'b0), .Q(
        \PR_add[5][17] ) );
  Flip_Flop \PR_add_reg[5][18]  ( .D(N526), .CLK(m1191), .R(1'b0), .Q(
        \PR_add[5][18] ) );
  Flip_Flop \PR_add_reg[5][19]  ( .D(N527), .CLK(m1191), .R(1'b0), .Q(
        \PR_add[5][19] ) );
  Flip_Flop \PR_add_reg[6][0]  ( .D(N528), .CLK(m1213), .R(1'b0), .Q(N248) );
  Flip_Flop \PR_add_reg[6][1]  ( .D(N529), .CLK(m1212), .R(1'b0), .Q(
        \PR_add[6][1] ) );
  Flip_Flop \PR_add_reg[6][2]  ( .D(N530), .CLK(m1210), .R(1'b0), .Q(
        \PR_add[6][2] ) );
  Flip_Flop \PR_add_reg[6][3]  ( .D(N531), .CLK(m1209), .R(1'b0), .Q(
        \PR_add[6][3] ) );
  Flip_Flop \PR_add_reg[6][4]  ( .D(N532), .CLK(m1208), .R(1'b0), .Q(
        \PR_add[6][4] ) );
  Flip_Flop \PR_add_reg[6][5]  ( .D(N533), .CLK(m1206), .R(1'b0), .Q(
        \PR_add[6][5] ) );
  Flip_Flop \PR_add_reg[6][6]  ( .D(N534), .CLK(m1205), .R(1'b0), .Q(
        \PR_add[6][6] ) );
  Flip_Flop \PR_add_reg[6][7]  ( .D(N535), .CLK(m1203), .R(1'b0), .Q(
        \PR_add[6][7] ) );
  Flip_Flop \PR_add_reg[6][8]  ( .D(N536), .CLK(m1202), .R(1'b0), .Q(
        \PR_add[6][8] ) );
  Flip_Flop \PR_add_reg[6][9]  ( .D(N537), .CLK(m1200), .R(1'b0), .Q(
        \PR_add[6][9] ) );
  Flip_Flop \PR_add_reg[6][10]  ( .D(N538), .CLK(m1198), .R(1'b0), .Q(
        \PR_add[6][10] ) );
  Flip_Flop \PR_add_reg[6][11]  ( .D(N539), .CLK(m1198), .R(1'b0), .Q(
        \PR_add[6][11] ) );
  Flip_Flop \PR_add_reg[6][12]  ( .D(N540), .CLK(m1196), .R(1'b0), .Q(
        \PR_add[6][12] ) );
  Flip_Flop \PR_add_reg[6][13]  ( .D(N541), .CLK(m1194), .R(1'b0), .Q(
        \PR_add[6][13] ) );
  Flip_Flop \PR_add_reg[6][14]  ( .D(N542), .CLK(m1193), .R(1'b0), .Q(
        \PR_add[6][14] ) );
  Flip_Flop \PR_add_reg[6][15]  ( .D(N543), .CLK(m1192), .R(1'b0), .Q(
        \PR_add[6][15] ) );
  Flip_Flop \PR_add_reg[6][16]  ( .D(N544), .CLK(m1191), .R(1'b0), .Q(
        \PR_add[6][16] ) );
  Flip_Flop \PR_add_reg[6][17]  ( .D(N545), .CLK(m1191), .R(1'b0), .Q(
        \PR_add[6][17] ) );
  Flip_Flop \PR_add_reg[6][18]  ( .D(N546), .CLK(m1191), .R(1'b0), .Q(
        \PR_add[6][18] ) );
  Flip_Flop \PR_add_reg[6][19]  ( .D(N547), .CLK(m1191), .R(1'b0), .Q(
        \PR_add[6][19] ) );
  Flip_Flop \PR_add_reg[7][0]  ( .D(N548), .CLK(m1213), .R(1'b0), .Q(N268) );
  Flip_Flop \PR_add_reg[7][1]  ( .D(N549), .CLK(m1212), .R(1'b0), .Q(N269) );
  Flip_Flop \PR_add_reg[7][2]  ( .D(N550), .CLK(m1210), .R(1'b0), .Q(
        \PR_add[7][2] ) );
  Flip_Flop \PR_add_reg[7][3]  ( .D(N551), .CLK(m1209), .R(1'b0), .Q(
        \PR_add[7][3] ) );
  Flip_Flop \PR_add_reg[7][4]  ( .D(N552), .CLK(m1207), .R(1'b0), .Q(
        \PR_add[7][4] ) );
  Flip_Flop \PR_add_reg[7][5]  ( .D(N553), .CLK(m1206), .R(1'b0), .Q(
        \PR_add[7][5] ) );
  Flip_Flop \PR_add_reg[7][6]  ( .D(N554), .CLK(m1205), .R(1'b0), .Q(
        \PR_add[7][6] ) );
  Flip_Flop \PR_add_reg[7][7]  ( .D(N555), .CLK(m1203), .R(1'b0), .Q(
        \PR_add[7][7] ) );
  Flip_Flop \PR_add_reg[7][8]  ( .D(N556), .CLK(m1202), .R(1'b0), .Q(
        \PR_add[7][8] ) );
  Flip_Flop \PR_add_reg[7][9]  ( .D(N557), .CLK(m1200), .R(1'b0), .Q(
        \PR_add[7][9] ) );
  Flip_Flop \PR_add_reg[7][10]  ( .D(N558), .CLK(m1198), .R(1'b0), .Q(
        \PR_add[7][10] ) );
  Flip_Flop \PR_add_reg[7][11]  ( .D(N559), .CLK(m1198), .R(1'b0), .Q(
        \PR_add[7][11] ) );
  Flip_Flop \PR_add_reg[7][12]  ( .D(N560), .CLK(m1196), .R(1'b0), .Q(
        \PR_add[7][12] ) );
  Flip_Flop \PR_add_reg[7][13]  ( .D(N561), .CLK(m1194), .R(1'b0), .Q(
        \PR_add[7][13] ) );
  Flip_Flop \PR_add_reg[7][14]  ( .D(N562), .CLK(m1193), .R(1'b0), .Q(
        \PR_add[7][14] ) );
  Flip_Flop \PR_add_reg[7][15]  ( .D(N563), .CLK(m1192), .R(1'b0), .Q(
        \PR_add[7][15] ) );
  Flip_Flop \PR_add_reg[7][16]  ( .D(N564), .CLK(m1190), .R(1'b0), .Q(
        \PR_add[7][16] ) );
  Flip_Flop \PR_add_reg[7][17]  ( .D(N565), .CLK(m1190), .R(1'b0), .Q(
        \PR_add[7][17] ) );
  Flip_Flop \PR_add_reg[7][18]  ( .D(N566), .CLK(m1190), .R(1'b0), .Q(
        \PR_add[7][18] ) );
  Flip_Flop \PR_add_reg[7][19]  ( .D(N567), .CLK(m1190), .R(1'b0), .Q(
        \PR_add[7][19] ) );
  Flip_Flop \PR_add_reg[8][0]  ( .D(N568), .CLK(m1213), .R(1'b0), .Q(
        \PR_add[8][0] ) );
  Flip_Flop \PR_add_reg[8][1]  ( .D(N569), .CLK(m1212), .R(1'b0), .Q(
        \PR_add[8][1] ) );
  Flip_Flop \PR_add_reg[8][2]  ( .D(N570), .CLK(m1210), .R(1'b0), .Q(
        \PR_add[8][2] ) );
  Flip_Flop \PR_add_reg[8][3]  ( .D(N571), .CLK(m1209), .R(1'b0), .Q(
        \PR_add[8][3] ) );
  Flip_Flop \PR_add_reg[8][4]  ( .D(N572), .CLK(m1207), .R(1'b0), .Q(
        \PR_add[8][4] ) );
  Flip_Flop \PR_add_reg[8][5]  ( .D(N573), .CLK(m1206), .R(1'b0), .Q(
        \PR_add[8][5] ) );
  Flip_Flop \PR_add_reg[8][6]  ( .D(N574), .CLK(m1205), .R(1'b0), .Q(
        \PR_add[8][6] ) );
  Flip_Flop \PR_add_reg[8][7]  ( .D(N575), .CLK(m1203), .R(1'b0), .Q(
        \PR_add[8][7] ) );
  Flip_Flop \PR_add_reg[8][8]  ( .D(N576), .CLK(m1202), .R(1'b0), .Q(
        \PR_add[8][8] ) );
  Flip_Flop \PR_add_reg[8][9]  ( .D(N577), .CLK(m1200), .R(1'b0), .Q(
        \PR_add[8][9] ) );
  Flip_Flop \PR_add_reg[8][10]  ( .D(N578), .CLK(m1197), .R(1'b0), .Q(
        \PR_add[8][10] ) );
  Flip_Flop \PR_add_reg[8][11]  ( .D(N579), .CLK(m1197), .R(1'b0), .Q(
        \PR_add[8][11] ) );
  Flip_Flop \PR_add_reg[8][12]  ( .D(N580), .CLK(m1196), .R(1'b0), .Q(
        \PR_add[8][12] ) );
  Flip_Flop \PR_add_reg[8][13]  ( .D(N581), .CLK(m1194), .R(1'b0), .Q(
        \PR_add[8][13] ) );
  Flip_Flop \PR_add_reg[8][14]  ( .D(N582), .CLK(m1193), .R(1'b0), .Q(
        \PR_add[8][14] ) );
  Flip_Flop \PR_add_reg[8][15]  ( .D(N583), .CLK(m1192), .R(1'b0), .Q(
        \PR_add[8][15] ) );
  Flip_Flop \PR_add_reg[8][16]  ( .D(N584), .CLK(m1190), .R(1'b0), .Q(
        \PR_add[8][16] ) );
  Flip_Flop \PR_add_reg[8][17]  ( .D(N585), .CLK(m1190), .R(1'b0), .Q(
        \PR_add[8][17] ) );
  Flip_Flop \PR_add_reg[8][18]  ( .D(N586), .CLK(m1190), .R(1'b0), .Q(
        \PR_add[8][18] ) );
  Flip_Flop \PR_add_reg[8][19]  ( .D(N587), .CLK(m1190), .R(1'b0), .Q(
        \PR_add[8][19] ) );
  Flip_Flop \PR_add_reg[9][0]  ( .D(N588), .CLK(m1213), .R(1'b0), .Q(N308) );
  Flip_Flop \PR_add_reg[9][1]  ( .D(N589), .CLK(m1212), .R(1'b0), .Q(N309) );
  Flip_Flop \PR_add_reg[9][2]  ( .D(N590), .CLK(m1210), .R(1'b0), .Q(N310) );
  Flip_Flop \PR_add_reg[9][3]  ( .D(N591), .CLK(m1209), .R(1'b0), .Q(
        \PR_add[9][3] ) );
  Flip_Flop \PR_add_reg[9][4]  ( .D(N592), .CLK(m1207), .R(1'b0), .Q(
        \PR_add[9][4] ) );
  Flip_Flop \PR_add_reg[9][5]  ( .D(N593), .CLK(m1206), .R(1'b0), .Q(
        \PR_add[9][5] ) );
  Flip_Flop \PR_add_reg[9][6]  ( .D(N594), .CLK(m1204), .R(1'b0), .Q(
        \PR_add[9][6] ) );
  Flip_Flop \PR_add_reg[9][7]  ( .D(N595), .CLK(m1203), .R(1'b0), .Q(
        \PR_add[9][7] ) );
  Flip_Flop \PR_add_reg[9][8]  ( .D(N596), .CLK(m1202), .R(1'b0), .Q(
        \PR_add[9][8] ) );
  Flip_Flop \PR_add_reg[9][9]  ( .D(N597), .CLK(m1200), .R(1'b0), .Q(
        \PR_add[9][9] ) );
  Flip_Flop \PR_add_reg[9][10]  ( .D(N598), .CLK(m1197), .R(1'b0), .Q(
        \PR_add[9][10] ) );
  Flip_Flop \PR_add_reg[9][11]  ( .D(N599), .CLK(m1197), .R(1'b0), .Q(
        \PR_add[9][11] ) );
  Flip_Flop \PR_add_reg[9][12]  ( .D(N600), .CLK(m1196), .R(1'b0), .Q(
        \PR_add[9][12] ) );
  Flip_Flop \PR_add_reg[9][13]  ( .D(N601), .CLK(m1194), .R(1'b0), .Q(
        \PR_add[9][13] ) );
  Flip_Flop \PR_add_reg[9][14]  ( .D(N602), .CLK(m1193), .R(1'b0), .Q(
        \PR_add[9][14] ) );
  Flip_Flop \PR_add_reg[9][15]  ( .D(N603), .CLK(m1192), .R(1'b0), .Q(
        \PR_add[9][15] ) );
  Flip_Flop \PR_add_reg[9][16]  ( .D(N604), .CLK(m1190), .R(1'b0), .Q(
        \PR_add[9][16] ) );
  Flip_Flop \PR_add_reg[9][17]  ( .D(N605), .CLK(m1190), .R(1'b0), .Q(
        \PR_add[9][17] ) );
  Flip_Flop \PR_add_reg[9][18]  ( .D(N606), .CLK(m1190), .R(1'b0), .Q(
        \PR_add[9][18] ) );
  Flip_Flop \PR_add_reg[9][19]  ( .D(N607), .CLK(m1190), .R(1'b0), .Q(
        \PR_add[9][19] ) );
  Flip_Flop \PR_add_reg[10][0]  ( .D(N608), .CLK(m1213), .R(1'b0), .Q(
        \PR_add[10][0] ) );
  Flip_Flop \PR_add_reg[10][1]  ( .D(N609), .CLK(m1211), .R(1'b0), .Q(
        \PR_add[10][1] ) );
  Flip_Flop \PR_add_reg[10][2]  ( .D(N610), .CLK(m1210), .R(1'b0), .Q(
        \PR_add[10][2] ) );
  Flip_Flop \PR_add_reg[10][3]  ( .D(N611), .CLK(m1209), .R(1'b0), .Q(
        \PR_add[10][3] ) );
  Flip_Flop \PR_add_reg[10][4]  ( .D(N612), .CLK(m1207), .R(1'b0), .Q(
        \PR_add[10][4] ) );
  Flip_Flop \PR_add_reg[10][5]  ( .D(N613), .CLK(m1206), .R(1'b0), .Q(
        \PR_add[10][5] ) );
  Flip_Flop \PR_add_reg[10][6]  ( .D(N614), .CLK(m1204), .R(1'b0), .Q(
        \PR_add[10][6] ) );
  Flip_Flop \PR_add_reg[10][7]  ( .D(N615), .CLK(m1203), .R(1'b0), .Q(
        \PR_add[10][7] ) );
  Flip_Flop \PR_add_reg[10][8]  ( .D(N616), .CLK(m1202), .R(1'b0), .Q(
        \PR_add[10][8] ) );
  Flip_Flop \PR_add_reg[10][9]  ( .D(N617), .CLK(m1200), .R(1'b0), .Q(
        \PR_add[10][9] ) );
  Flip_Flop \PR_add_reg[10][10]  ( .D(N618), .CLK(m1197), .R(1'b0), .Q(
        \PR_add[10][10] ) );
  Flip_Flop \PR_add_reg[10][11]  ( .D(N619), .CLK(m1197), .R(1'b0), .Q(
        \PR_add[10][11] ) );
  Flip_Flop \PR_add_reg[10][12]  ( .D(N620), .CLK(m1196), .R(1'b0), .Q(
        \PR_add[10][12] ) );
  Flip_Flop \PR_add_reg[10][13]  ( .D(N621), .CLK(m1194), .R(1'b0), .Q(
        \PR_add[10][13] ) );
  Flip_Flop \PR_add_reg[10][14]  ( .D(N622), .CLK(m1193), .R(1'b0), .Q(
        \PR_add[10][14] ) );
  Flip_Flop \PR_add_reg[10][15]  ( .D(N623), .CLK(m1192), .R(1'b0), .Q(
        \PR_add[10][15] ) );
  Flip_Flop \PR_add_reg[10][16]  ( .D(N624), .CLK(m1189), .R(1'b0), .Q(
        \PR_add[10][16] ) );
  Flip_Flop \PR_add_reg[10][17]  ( .D(N625), .CLK(m1189), .R(1'b0), .Q(
        \PR_add[10][17] ) );
  Flip_Flop \PR_add_reg[10][18]  ( .D(N626), .CLK(m1189), .R(1'b0), .Q(
        \PR_add[10][18] ) );
  Flip_Flop \PR_add_reg[10][19]  ( .D(N627), .CLK(m1189), .R(1'b0), .Q(
        \PR_add[10][19] ) );
  Flip_Flop \PR_add_reg[11][0]  ( .D(N628), .CLK(m1213), .R(1'b0), .Q(N348) );
  Flip_Flop \PR_add_reg[11][1]  ( .D(N629), .CLK(m1211), .R(1'b0), .Q(
        \PR_add[11][1] ) );
  Flip_Flop \PR_add_reg[11][2]  ( .D(N630), .CLK(m1210), .R(1'b0), .Q(
        \PR_add[11][2] ) );
  Flip_Flop \PR_add_reg[11][3]  ( .D(N631), .CLK(m1209), .R(1'b0), .Q(
        \PR_add[11][3] ) );
  Flip_Flop \PR_add_reg[11][4]  ( .D(N632), .CLK(m1207), .R(1'b0), .Q(
        \PR_add[11][4] ) );
  Flip_Flop \PR_add_reg[11][5]  ( .D(N633), .CLK(m1206), .R(1'b0), .Q(
        \PR_add[11][5] ) );
  Flip_Flop \PR_add_reg[11][6]  ( .D(N634), .CLK(m1204), .R(1'b0), .Q(
        \PR_add[11][6] ) );
  Flip_Flop \PR_add_reg[11][7]  ( .D(N635), .CLK(m1203), .R(1'b0), .Q(
        \PR_add[11][7] ) );
  Flip_Flop \PR_add_reg[11][8]  ( .D(N636), .CLK(m1201), .R(1'b0), .Q(
        \PR_add[11][8] ) );
  Flip_Flop \PR_add_reg[11][9]  ( .D(N637), .CLK(m1200), .R(1'b0), .Q(
        \PR_add[11][9] ) );
  Flip_Flop \PR_add_reg[11][10]  ( .D(N638), .CLK(m1197), .R(1'b0), .Q(
        \PR_add[11][10] ) );
  Flip_Flop \PR_add_reg[11][11]  ( .D(N639), .CLK(m1197), .R(1'b0), .Q(
        \PR_add[11][11] ) );
  Flip_Flop \PR_add_reg[11][12]  ( .D(N640), .CLK(m1195), .R(1'b0), .Q(
        \PR_add[11][12] ) );
  Flip_Flop \PR_add_reg[11][13]  ( .D(N641), .CLK(m1194), .R(1'b0), .Q(
        \PR_add[11][13] ) );
  Flip_Flop \PR_add_reg[11][14]  ( .D(N642), .CLK(m1192), .R(1'b0), .Q(
        \PR_add[11][14] ) );
  Flip_Flop \PR_add_reg[11][15]  ( .D(N643), .CLK(m1192), .R(1'b0), .Q(
        \PR_add[11][15] ) );
  Flip_Flop \PR_add_reg[11][16]  ( .D(N644), .CLK(m1189), .R(1'b0), .Q(
        \PR_add[11][16] ) );
  Flip_Flop \PR_add_reg[11][17]  ( .D(N645), .CLK(m1189), .R(1'b0), .Q(
        \PR_add[11][17] ) );
  Flip_Flop \PR_add_reg[11][18]  ( .D(N646), .CLK(m1189), .R(1'b0), .Q(
        \PR_add[11][18] ) );
  Flip_Flop \PR_add_reg[11][19]  ( .D(N647), .CLK(m1189), .R(1'b0), .Q(
        \PR_add[11][19] ) );
  Flip_Flop \PR_add_reg[12][0]  ( .D(N648), .CLK(m1213), .R(1'b0), .Q(N368) );
  Flip_Flop \PR_add_reg[12][1]  ( .D(N649), .CLK(m1211), .R(1'b0), .Q(N369) );
  Flip_Flop \PR_add_reg[12][2]  ( .D(N650), .CLK(m1210), .R(1'b0), .Q(
        \PR_add[12][2] ) );
  Flip_Flop \PR_add_reg[12][3]  ( .D(N651), .CLK(m1208), .R(1'b0), .Q(
        \PR_add[12][3] ) );
  Flip_Flop \PR_add_reg[12][4]  ( .D(N652), .CLK(m1207), .R(1'b0), .Q(
        \PR_add[12][4] ) );
  Flip_Flop \PR_add_reg[12][5]  ( .D(N653), .CLK(m1206), .R(1'b0), .Q(
        \PR_add[12][5] ) );
  Flip_Flop \PR_add_reg[12][6]  ( .D(N654), .CLK(m1204), .R(1'b0), .Q(
        \PR_add[12][6] ) );
  Flip_Flop \PR_add_reg[12][7]  ( .D(N655), .CLK(m1203), .R(1'b0), .Q(
        \PR_add[12][7] ) );
  Flip_Flop \PR_add_reg[12][8]  ( .D(N656), .CLK(m1201), .R(1'b0), .Q(
        \PR_add[12][8] ) );
  Flip_Flop \PR_add_reg[12][9]  ( .D(N657), .CLK(m1200), .R(1'b0), .Q(
        \PR_add[12][9] ) );
  Flip_Flop \PR_add_reg[12][10]  ( .D(N658), .CLK(m1197), .R(1'b0), .Q(
        \PR_add[12][10] ) );
  Flip_Flop \PR_add_reg[12][11]  ( .D(N659), .CLK(m1197), .R(1'b0), .Q(
        \PR_add[12][11] ) );
  Flip_Flop \PR_add_reg[12][12]  ( .D(N660), .CLK(m1195), .R(1'b0), .Q(
        \PR_add[12][12] ) );
  Flip_Flop \PR_add_reg[12][13]  ( .D(N661), .CLK(m1194), .R(1'b0), .Q(
        \PR_add[12][13] ) );
  Flip_Flop \PR_add_reg[12][14]  ( .D(N662), .CLK(m1192), .R(1'b0), .Q(
        \PR_add[12][14] ) );
  Flip_Flop \PR_add_reg[12][15]  ( .D(N663), .CLK(m1191), .R(1'b0), .Q(
        \PR_add[12][15] ) );
  Flip_Flop \PR_add_reg[12][16]  ( .D(N664), .CLK(m1189), .R(1'b0), .Q(
        \PR_add[12][16] ) );
  Flip_Flop \PR_add_reg[12][17]  ( .D(N665), .CLK(m1189), .R(1'b0), .Q(
        \PR_add[12][17] ) );
  Flip_Flop \PR_add_reg[12][18]  ( .D(N666), .CLK(m1189), .R(1'b0), .Q(
        \PR_add[12][18] ) );
  Flip_Flop \PR_add_reg[12][19]  ( .D(N667), .CLK(m1189), .R(1'b0), .Q(
        \PR_add[12][19] ) );
  Flip_Flop \PR_add_reg[13][0]  ( .D(N668), .CLK(m1213), .R(1'b0), .Q(
        \PR_add[13][0] ) );
  Flip_Flop \acc_reg[0]  ( .D(N953), .CLK(m1213), .R(1'b0), .Q(acc[0]) );
  Flip_Flop \Data_out_reg[0]  ( .D(N388), .CLK(m1212), .R(1'b0), .Q(
        Data_out[0]) );
  Flip_Flop \PR_add_reg[13][1]  ( .D(N669), .CLK(m1211), .R(1'b0), .Q(
        \PR_add[13][1] ) );
  Flip_Flop \acc_reg[1]  ( .D(N954), .CLK(m1211), .R(1'b0), .Q(acc[1]) );
  Flip_Flop \Data_out_reg[1]  ( .D(N389), .CLK(m1211), .R(1'b0), .Q(
        Data_out[1]) );
  Flip_Flop \PR_add_reg[13][2]  ( .D(N670), .CLK(m1210), .R(1'b0), .Q(
        \PR_add[13][2] ) );
  Flip_Flop \acc_reg[2]  ( .D(N955), .CLK(m1210), .R(1'b0), .Q(acc[2]) );
  Flip_Flop \Data_out_reg[2]  ( .D(N390), .CLK(m1210), .R(1'b0), .Q(
        Data_out[2]) );
  Flip_Flop \PR_add_reg[13][3]  ( .D(N671), .CLK(m1208), .R(1'b0), .Q(
        \PR_add[13][3] ) );
  Flip_Flop \acc_reg[3]  ( .D(N956), .CLK(m1208), .R(1'b0), .Q(acc[3]) );
  Flip_Flop \Data_out_reg[3]  ( .D(N391), .CLK(m1208), .R(1'b0), .Q(
        Data_out[3]) );
  Flip_Flop \PR_add_reg[13][4]  ( .D(N672), .CLK(m1207), .R(1'b0), .Q(
        \PR_add[13][4] ) );
  Flip_Flop \acc_reg[4]  ( .D(N957), .CLK(m1207), .R(1'b0), .Q(acc[4]) );
  Flip_Flop \Data_out_reg[4]  ( .D(N392), .CLK(m1207), .R(1'b0), .Q(
        Data_out[4]) );
  Flip_Flop \PR_add_reg[13][5]  ( .D(N673), .CLK(m1206), .R(1'b0), .Q(
        \PR_add[13][5] ) );
  Flip_Flop \acc_reg[5]  ( .D(N958), .CLK(m1205), .R(1'b0), .Q(acc[5]) );
  Flip_Flop \Data_out_reg[5]  ( .D(N393), .CLK(m1205), .R(1'b0), .Q(
        Data_out[5]) );
  Flip_Flop \PR_add_reg[13][6]  ( .D(N674), .CLK(m1204), .R(1'b0), .Q(
        \PR_add[13][6] ) );
  Flip_Flop \acc_reg[6]  ( .D(N959), .CLK(m1204), .R(1'b0), .Q(acc[6]) );
  Flip_Flop \Data_out_reg[6]  ( .D(N394), .CLK(m1204), .R(1'b0), .Q(
        Data_out[6]) );
  Flip_Flop \PR_add_reg[13][7]  ( .D(N675), .CLK(m1203), .R(1'b0), .Q(
        \PR_add[13][7] ) );
  Flip_Flop \acc_reg[7]  ( .D(N960), .CLK(m1203), .R(1'b0), .Q(acc[7]) );
  Flip_Flop \Data_out_reg[7]  ( .D(N395), .CLK(m1203), .R(1'b0), .Q(
        Data_out[7]) );
  Flip_Flop \PR_add_reg[13][8]  ( .D(N676), .CLK(m1201), .R(1'b0), .Q(
        \PR_add[13][8] ) );
  Flip_Flop \acc_reg[8]  ( .D(N961), .CLK(m1201), .R(1'b0), .Q(acc[8]) );
  Flip_Flop \Data_out_reg[8]  ( .D(N396), .CLK(m1201), .R(1'b0), .Q(
        Data_out[8]) );
  Flip_Flop \PR_add_reg[13][9]  ( .D(N677), .CLK(m1200), .R(1'b0), .Q(
        \PR_add[13][9] ) );
  Flip_Flop \acc_reg[9]  ( .D(N962), .CLK(m1200), .R(1'b0), .Q(acc[9]) );
  Flip_Flop \Data_out_reg[9]  ( .D(N397), .CLK(m1200), .R(1'b0), .Q(
        Data_out[9]) );
  Flip_Flop \PR_add_reg[13][10]  ( .D(N678), .CLK(m1196), .R(1'b0), .Q(
        \PR_add[13][10] ) );
  Flip_Flop \acc_reg[10]  ( .D(N963), .CLK(m1196), .R(1'b0), .Q(acc[10]) );
  Flip_Flop \Data_out_reg[10]  ( .D(N398), .CLK(m1196), .R(1'b0), .Q(
        Data_out[10]) );
  Flip_Flop \PR_add_reg[13][11]  ( .D(N679), .CLK(m1197), .R(1'b0), .Q(
        \PR_add[13][11] ) );
  Flip_Flop \acc_reg[11]  ( .D(N964), .CLK(m1197), .R(1'b0), .Q(acc[11]) );
  Flip_Flop \Data_out_reg[11]  ( .D(N399), .CLK(m1196), .R(1'b0), .Q(
        Data_out[11]) );
  Flip_Flop \PR_add_reg[13][12]  ( .D(N680), .CLK(m1195), .R(1'b0), .Q(
        \PR_add[13][12] ) );
  Flip_Flop \acc_reg[12]  ( .D(N965), .CLK(m1195), .R(1'b0), .Q(acc[12]) );
  Flip_Flop \Data_out_reg[12]  ( .D(N400), .CLK(m1195), .R(1'b0), .Q(
        Data_out[12]) );
  Flip_Flop \PR_add_reg[13][13]  ( .D(N681), .CLK(m1194), .R(1'b0), .Q(
        \PR_add[13][13] ) );
  Flip_Flop \acc_reg[13]  ( .D(N966), .CLK(m1194), .R(1'b0), .Q(acc[13]) );
  Flip_Flop \Data_out_reg[13]  ( .D(N401), .CLK(m1194), .R(1'b0), .Q(
        Data_out[13]) );
  Flip_Flop \PR_add_reg[13][14]  ( .D(N682), .CLK(m1192), .R(1'b0), .Q(
        \PR_add[13][14] ) );
  Flip_Flop \acc_reg[14]  ( .D(N967), .CLK(m1192), .R(1'b0), .Q(acc[14]) );
  Flip_Flop \Data_out_reg[14]  ( .D(N402), .CLK(m1192), .R(1'b0), .Q(
        Data_out[14]) );
  Flip_Flop \PR_add_reg[13][15]  ( .D(N683), .CLK(m1191), .R(1'b0), .Q(
        \PR_add[13][15] ) );
  Flip_Flop \acc_reg[15]  ( .D(N968), .CLK(m1191), .R(1'b0), .Q(acc[15]) );
  Flip_Flop \Data_out_reg[15]  ( .D(N403), .CLK(m1191), .R(1'b0), .Q(
        Data_out[15]) );
  Flip_Flop \PR_add_reg[13][16]  ( .D(N684), .CLK(m1188), .R(1'b0), .Q(
        \PR_add[13][16] ) );
  Flip_Flop \acc_reg[16]  ( .D(N969), .CLK(m1188), .R(1'b0), .Q(acc[16]) );
  Flip_Flop \Data_out_reg[16]  ( .D(N404), .CLK(m1188), .R(1'b0), .Q(
        Data_out[16]) );
  Flip_Flop \PR_add_reg[13][17]  ( .D(N685), .CLK(m1188), .R(1'b0), .Q(
        \PR_add[13][17] ) );
  Flip_Flop \acc_reg[17]  ( .D(N970), .CLK(m1188), .R(1'b0), .Q(acc[17]) );
  Flip_Flop \Data_out_reg[17]  ( .D(N405), .CLK(m1188), .R(1'b0), .Q(
        Data_out[17]) );
  Flip_Flop \PR_add_reg[13][18]  ( .D(N686), .CLK(m1188), .R(1'b0), .Q(
        \PR_add[13][18] ) );
  Flip_Flop \acc_reg[18]  ( .D(N971), .CLK(m1188), .R(1'b0), .Q(acc[18]) );
  Flip_Flop \Data_out_reg[18]  ( .D(N406), .CLK(m1188), .R(1'b0), .Q(
        Data_out[18]) );
  Flip_Flop \PR_add_reg[13][19]  ( .D(N687), .CLK(m1188), .R(1'b0), .Q(
        \PR_add[13][19] ) );
  Flip_Flop \acc_reg[19]  ( .D(N972), .CLK(m1188), .R(1'b0), .Q(acc[19]) );
  Flip_Flop \Data_out_reg[19]  ( .D(N407), .CLK(m1188), .R(1'b0), .Q(
        Data_out[19]) );
  INV U610 ( .IN(clock), .OUT(m631) );
  NOR2 U759 ( .A(m1252), .B(m633), .OUT(N972) );
  INV U760 ( .IN(\PR_add[13][19] ), .OUT(m633) );
  NOR2 U761 ( .A(m1252), .B(m634), .OUT(N971) );
  INV U762 ( .IN(\PR_add[13][18] ), .OUT(m634) );
  NOR2 U763 ( .A(m1252), .B(m635), .OUT(N970) );
  INV U764 ( .IN(\PR_add[13][17] ), .OUT(m635) );
  NOR2 U765 ( .A(m1252), .B(m636), .OUT(N969) );
  INV U766 ( .IN(\PR_add[13][16] ), .OUT(m636) );
  NOR2 U767 ( .A(m1252), .B(m637), .OUT(N968) );
  INV U768 ( .IN(\PR_add[13][15] ), .OUT(m637) );
  NOR2 U769 ( .A(m1252), .B(m638), .OUT(N967) );
  INV U770 ( .IN(\PR_add[13][14] ), .OUT(m638) );
  NOR2 U771 ( .A(m1252), .B(m639), .OUT(N966) );
  INV U772 ( .IN(\PR_add[13][13] ), .OUT(m639) );
  NOR2 U773 ( .A(m1252), .B(m640), .OUT(N965) );
  INV U774 ( .IN(\PR_add[13][12] ), .OUT(m640) );
  NOR2 U775 ( .A(m1252), .B(m641), .OUT(N964) );
  INV U776 ( .IN(\PR_add[13][11] ), .OUT(m641) );
  NOR2 U777 ( .A(m1252), .B(m642), .OUT(N963) );
  INV U778 ( .IN(\PR_add[13][10] ), .OUT(m642) );
  NOR2 U779 ( .A(m1252), .B(m643), .OUT(N962) );
  INV U780 ( .IN(\PR_add[13][9] ), .OUT(m643) );
  NOR2 U781 ( .A(m1252), .B(m644), .OUT(N961) );
  INV U782 ( .IN(\PR_add[13][8] ), .OUT(m644) );
  NOR2 U783 ( .A(m1252), .B(m645), .OUT(N960) );
  INV U784 ( .IN(\PR_add[13][7] ), .OUT(m645) );
  NOR2 U785 ( .A(m1253), .B(m646), .OUT(N959) );
  INV U786 ( .IN(\PR_add[13][6] ), .OUT(m646) );
  NOR2 U787 ( .A(m1253), .B(m647), .OUT(N958) );
  INV U788 ( .IN(\PR_add[13][5] ), .OUT(m647) );
  NOR2 U789 ( .A(m1253), .B(m648), .OUT(N957) );
  INV U790 ( .IN(\PR_add[13][4] ), .OUT(m648) );
  NOR2 U791 ( .A(m1253), .B(m649), .OUT(N956) );
  INV U792 ( .IN(\PR_add[13][3] ), .OUT(m649) );
  NOR2 U793 ( .A(m1253), .B(m650), .OUT(N955) );
  INV U794 ( .IN(\PR_add[13][2] ), .OUT(m650) );
  NOR2 U795 ( .A(m1253), .B(m651), .OUT(N954) );
  INV U796 ( .IN(\PR_add[13][1] ), .OUT(m651) );
  NOR2 U797 ( .A(m1253), .B(m652), .OUT(N953) );
  INV U798 ( .IN(\PR_add[13][0] ), .OUT(m652) );
  NOR2 U799 ( .A(m1253), .B(m653), .OUT(N952) );
  INV U800 ( .IN(\Samples[13][7] ), .OUT(m653) );
  NOR2 U801 ( .A(m1253), .B(m654), .OUT(N951) );
  INV U802 ( .IN(\Samples[13][6] ), .OUT(m654) );
  NOR2 U803 ( .A(m1253), .B(m655), .OUT(N950) );
  INV U804 ( .IN(\Samples[13][5] ), .OUT(m655) );
  NOR2 U805 ( .A(m1253), .B(m656), .OUT(N949) );
  INV U806 ( .IN(\Samples[13][4] ), .OUT(m656) );
  NOR2 U807 ( .A(m1253), .B(m657), .OUT(N948) );
  INV U808 ( .IN(\Samples[13][3] ), .OUT(m657) );
  NOR2 U809 ( .A(m1253), .B(m658), .OUT(N947) );
  INV U810 ( .IN(\Samples[13][2] ), .OUT(m658) );
  NOR2 U811 ( .A(m1254), .B(m659), .OUT(N946) );
  INV U812 ( .IN(\Samples[13][1] ), .OUT(m659) );
  NOR2 U813 ( .A(m1254), .B(m660), .OUT(N945) );
  INV U814 ( .IN(\Samples[13][0] ), .OUT(m660) );
  NOR2 U815 ( .A(m1254), .B(m661), .OUT(N944) );
  INV U816 ( .IN(N107), .OUT(m661) );
  NOR2 U817 ( .A(m1254), .B(m662), .OUT(N943) );
  INV U818 ( .IN(N106), .OUT(m662) );
  NOR2 U819 ( .A(m1254), .B(m663), .OUT(N942) );
  INV U820 ( .IN(N105), .OUT(m663) );
  NOR2 U821 ( .A(m1254), .B(m664), .OUT(N941) );
  INV U822 ( .IN(N104), .OUT(m664) );
  NOR2 U823 ( .A(m1254), .B(m665), .OUT(N940) );
  INV U824 ( .IN(N103), .OUT(m665) );
  NOR2 U825 ( .A(m1254), .B(m666), .OUT(N939) );
  INV U826 ( .IN(N102), .OUT(m666) );
  NOR2 U827 ( .A(m1254), .B(m667), .OUT(N938) );
  INV U828 ( .IN(N101), .OUT(m667) );
  NOR2 U829 ( .A(m1254), .B(m668), .OUT(N937) );
  INV U830 ( .IN(N100), .OUT(m668) );
  NOR2 U831 ( .A(m1254), .B(m669), .OUT(N936) );
  INV U832 ( .IN(N99), .OUT(m669) );
  NOR2 U833 ( .A(m1254), .B(m670), .OUT(N935) );
  INV U834 ( .IN(N98), .OUT(m670) );
  NOR2 U839 ( .A(m1254), .B(m673), .OUT(N932) );
  INV U840 ( .IN(N95), .OUT(m673) );
  NOR2 U841 ( .A(m1255), .B(m674), .OUT(N931) );
  INV U842 ( .IN(N94), .OUT(m674) );
  NOR2 U843 ( .A(m1255), .B(m675), .OUT(N930) );
  INV U844 ( .IN(N93), .OUT(m675) );
  NOR2 U845 ( .A(m1255), .B(m676), .OUT(N929) );
  INV U846 ( .IN(N92), .OUT(m676) );
  NOR2 U847 ( .A(m1255), .B(m677), .OUT(N928) );
  INV U848 ( .IN(N91), .OUT(m677) );
  NOR2 U849 ( .A(m1255), .B(m678), .OUT(N927) );
  INV U850 ( .IN(N90), .OUT(m678) );
  NOR2 U851 ( .A(m1255), .B(m679), .OUT(N926) );
  INV U852 ( .IN(N89), .OUT(m679) );
  NOR2 U853 ( .A(m1255), .B(m680), .OUT(N925) );
  INV U854 ( .IN(N88), .OUT(m680) );
  NOR2 U855 ( .A(m1255), .B(m681), .OUT(N924) );
  INV U856 ( .IN(N87), .OUT(m681) );
  NOR2 U857 ( .A(m1255), .B(m682), .OUT(N923) );
  INV U858 ( .IN(N86), .OUT(m682) );
  NOR2 U859 ( .A(m1255), .B(m683), .OUT(N922) );
  INV U860 ( .IN(N85), .OUT(m683) );
  NOR2 U861 ( .A(m1255), .B(m684), .OUT(N921) );
  INV U862 ( .IN(N84), .OUT(m684) );
  NOR2 U863 ( .A(m1255), .B(m685), .OUT(N912) );
  INV U864 ( .IN(N83), .OUT(m685) );
  NOR2 U865 ( .A(m1255), .B(m686), .OUT(N911) );
  INV U866 ( .IN(N82), .OUT(m686) );
  NOR2 U867 ( .A(m1256), .B(m687), .OUT(N910) );
  INV U868 ( .IN(N81), .OUT(m687) );
  NOR2 U869 ( .A(m1256), .B(m688), .OUT(N909) );
  INV U870 ( .IN(N80), .OUT(m688) );
  NOR2 U871 ( .A(m1256), .B(m689), .OUT(N908) );
  INV U872 ( .IN(N79), .OUT(m689) );
  NOR2 U873 ( .A(m1256), .B(m690), .OUT(N907) );
  INV U874 ( .IN(N78), .OUT(m690) );
  NOR2 U875 ( .A(m1256), .B(m691), .OUT(N906) );
  INV U876 ( .IN(N77), .OUT(m691) );
  NOR2 U877 ( .A(m1256), .B(m692), .OUT(N905) );
  INV U878 ( .IN(N76), .OUT(m692) );
  NOR2 U879 ( .A(m1256), .B(m693), .OUT(N904) );
  INV U880 ( .IN(N75), .OUT(m693) );
  NOR2 U881 ( .A(m1256), .B(m694), .OUT(N903) );
  INV U882 ( .IN(N74), .OUT(m694) );
  NOR2 U883 ( .A(m1256), .B(m695), .OUT(N902) );
  INV U884 ( .IN(N73), .OUT(m695) );
  NOR2 U885 ( .A(m1256), .B(m696), .OUT(N893) );
  INV U886 ( .IN(N72), .OUT(m696) );
  NOR2 U887 ( .A(m1256), .B(m697), .OUT(N892) );
  INV U888 ( .IN(N71), .OUT(m697) );
  NOR2 U889 ( .A(m1256), .B(m698), .OUT(N891) );
  INV U890 ( .IN(N70), .OUT(m698) );
  NOR2 U891 ( .A(m1256), .B(m699), .OUT(N890) );
  INV U892 ( .IN(N69), .OUT(m699) );
  NOR2 U893 ( .A(m1257), .B(m700), .OUT(N889) );
  INV U894 ( .IN(N68), .OUT(m700) );
  NOR2 U895 ( .A(m1257), .B(m701), .OUT(N888) );
  INV U896 ( .IN(N67), .OUT(m701) );
  NOR2 U897 ( .A(m1257), .B(m702), .OUT(N887) );
  INV U898 ( .IN(N66), .OUT(m702) );
  NOR2 U899 ( .A(m1257), .B(m703), .OUT(N886) );
  INV U900 ( .IN(N65), .OUT(m703) );
  NOR2 U901 ( .A(m1257), .B(m704), .OUT(N885) );
  INV U902 ( .IN(N64), .OUT(m704) );
  NOR2 U903 ( .A(m1257), .B(m705), .OUT(N884) );
  INV U904 ( .IN(N63), .OUT(m705) );
  NOR2 U909 ( .A(m1257), .B(m708), .OUT(N881) );
  INV U910 ( .IN(N60), .OUT(m708) );
  NOR2 U911 ( .A(m1257), .B(m709), .OUT(N880) );
  INV U912 ( .IN(N59), .OUT(m709) );
  NOR2 U913 ( .A(m1257), .B(m710), .OUT(N879) );
  INV U914 ( .IN(N58), .OUT(m710) );
  NOR2 U915 ( .A(m1257), .B(m711), .OUT(N878) );
  INV U916 ( .IN(N57), .OUT(m711) );
  NOR2 U917 ( .A(m1257), .B(m712), .OUT(N877) );
  INV U918 ( .IN(N56), .OUT(m712) );
  NOR2 U919 ( .A(m1257), .B(m713), .OUT(N876) );
  INV U920 ( .IN(N55), .OUT(m713) );
  NOR2 U921 ( .A(m1257), .B(m714), .OUT(N875) );
  INV U922 ( .IN(N54), .OUT(m714) );
  NOR2 U923 ( .A(m1258), .B(m715), .OUT(N874) );
  INV U924 ( .IN(N53), .OUT(m715) );
  NOR2 U925 ( .A(m1258), .B(m716), .OUT(N873) );
  INV U926 ( .IN(N52), .OUT(m716) );
  NOR2 U927 ( .A(m1258), .B(m717), .OUT(N872) );
  INV U928 ( .IN(N51), .OUT(m717) );
  NOR2 U929 ( .A(m1258), .B(m718), .OUT(N871) );
  INV U930 ( .IN(N50), .OUT(m718) );
  NOR2 U931 ( .A(m1258), .B(m719), .OUT(N870) );
  INV U932 ( .IN(N49), .OUT(m719) );
  NOR2 U933 ( .A(m1258), .B(m720), .OUT(N861) );
  INV U934 ( .IN(N48), .OUT(m720) );
  NOR2 U935 ( .A(m1258), .B(m721), .OUT(N860) );
  INV U936 ( .IN(N47), .OUT(m721) );
  NOR2 U937 ( .A(m1258), .B(m722), .OUT(N859) );
  INV U938 ( .IN(N46), .OUT(m722) );
  NOR2 U939 ( .A(m1258), .B(m723), .OUT(N858) );
  INV U940 ( .IN(N45), .OUT(m723) );
  NOR2 U941 ( .A(m1258), .B(m724), .OUT(N857) );
  INV U942 ( .IN(N44), .OUT(m724) );
  NOR2 U943 ( .A(m1258), .B(m725), .OUT(N856) );
  INV U944 ( .IN(N43), .OUT(m725) );
  NOR2 U945 ( .A(m1258), .B(m726), .OUT(N855) );
  INV U946 ( .IN(N42), .OUT(m726) );
  NOR2 U947 ( .A(m1258), .B(m727), .OUT(N854) );
  INV U948 ( .IN(N41), .OUT(m727) );
  NOR2 U949 ( .A(m1259), .B(m728), .OUT(N853) );
  INV U950 ( .IN(N40), .OUT(m728) );
  NOR2 U951 ( .A(m1259), .B(m729), .OUT(N852) );
  INV U952 ( .IN(N39), .OUT(m729) );
  NOR2 U953 ( .A(m1259), .B(m730), .OUT(N851) );
  INV U954 ( .IN(N38), .OUT(m730) );
  NOR2 U955 ( .A(m1259), .B(m731), .OUT(N842) );
  INV U956 ( .IN(N37), .OUT(m731) );
  NOR2 U957 ( .A(m1259), .B(m732), .OUT(N841) );
  INV U958 ( .IN(N36), .OUT(m732) );
  NOR2 U959 ( .A(m1259), .B(m733), .OUT(N840) );
  INV U960 ( .IN(N35), .OUT(m733) );
  NOR2 U961 ( .A(m1259), .B(m734), .OUT(N839) );
  INV U962 ( .IN(N34), .OUT(m734) );
  NOR2 U963 ( .A(m1259), .B(m735), .OUT(N838) );
  INV U964 ( .IN(N33), .OUT(m735) );
  NOR2 U965 ( .A(m1259), .B(m736), .OUT(N837) );
  INV U966 ( .IN(N32), .OUT(m736) );
  NOR2 U967 ( .A(m1259), .B(m737), .OUT(N836) );
  INV U968 ( .IN(N31), .OUT(m737) );
  NOR2 U969 ( .A(m1259), .B(m738), .OUT(N835) );
  INV U970 ( .IN(N30), .OUT(m738) );
  NOR2 U971 ( .A(m1259), .B(m739), .OUT(N834) );
  INV U972 ( .IN(N29), .OUT(m739) );
  NOR2 U973 ( .A(m1259), .B(m740), .OUT(N833) );
  INV U974 ( .IN(N28), .OUT(m740) );
  NOR2 U979 ( .A(m1260), .B(m743), .OUT(N830) );
  INV U980 ( .IN(N25), .OUT(m743) );
  NOR2 U981 ( .A(m1260), .B(m744), .OUT(N829) );
  INV U982 ( .IN(N24), .OUT(m744) );
  NOR2 U983 ( .A(m1260), .B(m745), .OUT(N828) );
  INV U984 ( .IN(N23), .OUT(m745) );
  NOR2 U985 ( .A(m1260), .B(m746), .OUT(N827) );
  INV U986 ( .IN(N22), .OUT(m746) );
  NOR2 U987 ( .A(m1260), .B(m747), .OUT(N826) );
  INV U988 ( .IN(N21), .OUT(m747) );
  NOR2 U989 ( .A(m1260), .B(m748), .OUT(N825) );
  INV U990 ( .IN(N20), .OUT(m748) );
  NOR2 U991 ( .A(m1260), .B(m749), .OUT(N824) );
  INV U992 ( .IN(N19), .OUT(m749) );
  NOR2 U993 ( .A(m1260), .B(m750), .OUT(N823) );
  INV U994 ( .IN(N18), .OUT(m750) );
  NOR2 U995 ( .A(m1260), .B(m751), .OUT(N822) );
  INV U996 ( .IN(N17), .OUT(m751) );
  NOR2 U997 ( .A(m1260), .B(m752), .OUT(N821) );
  INV U998 ( .IN(N16), .OUT(m752) );
  NOR2 U999 ( .A(m1260), .B(m753), .OUT(N820) );
  INV U1000 ( .IN(N15), .OUT(m753) );
  NOR2 U1001 ( .A(m1260), .B(m754), .OUT(N819) );
  INV U1002 ( .IN(N14), .OUT(m754) );
  NOR2 U1003 ( .A(m1260), .B(m755), .OUT(N810) );
  INV U1004 ( .IN(N13), .OUT(m755) );
  NOR2 U1005 ( .A(m1261), .B(m756), .OUT(N809) );
  INV U1006 ( .IN(N12), .OUT(m756) );
  NOR2 U1007 ( .A(m1261), .B(m757), .OUT(N808) );
  INV U1008 ( .IN(N11), .OUT(m757) );
  NOR2 U1009 ( .A(m1261), .B(m758), .OUT(N807) );
  INV U1010 ( .IN(N10), .OUT(m758) );
  NOR2 U1011 ( .A(m1261), .B(m759), .OUT(N806) );
  INV U1012 ( .IN(N9), .OUT(m759) );
  NOR2 U1013 ( .A(m1261), .B(m760), .OUT(N805) );
  INV U1014 ( .IN(N8), .OUT(m760) );
  NOR2 U1015 ( .A(m1261), .B(m761), .OUT(N804) );
  INV U1016 ( .IN(N7), .OUT(m761) );
  NOR2 U1017 ( .A(m1261), .B(m762), .OUT(N803) );
  INV U1018 ( .IN(N6), .OUT(m762) );
  NOR2 U1019 ( .A(m1261), .B(m763), .OUT(N802) );
  INV U1020 ( .IN(N5), .OUT(m763) );
  NOR2 U1021 ( .A(m1261), .B(m764), .OUT(N801) );
  INV U1022 ( .IN(N4), .OUT(m764) );
  NOR2 U1023 ( .A(m1261), .B(m765), .OUT(N800) );
  INV U1024 ( .IN(N3), .OUT(m765) );
  NOR2 U1025 ( .A(m1261), .B(m766), .OUT(N799) );
  INV U1026 ( .IN(\Samples[12][7] ), .OUT(m766) );
  NOR2 U1027 ( .A(m1261), .B(m767), .OUT(N798) );
  INV U1028 ( .IN(\Samples[12][6] ), .OUT(m767) );
  NOR2 U1029 ( .A(m1261), .B(m768), .OUT(N797) );
  INV U1030 ( .IN(\Samples[12][5] ), .OUT(m768) );
  NOR2 U1031 ( .A(m1262), .B(m769), .OUT(N796) );
  INV U1032 ( .IN(\Samples[12][4] ), .OUT(m769) );
  NOR2 U1033 ( .A(m1262), .B(m770), .OUT(N795) );
  INV U1034 ( .IN(\Samples[12][3] ), .OUT(m770) );
  NOR2 U1035 ( .A(m1262), .B(m771), .OUT(N794) );
  INV U1036 ( .IN(\Samples[12][2] ), .OUT(m771) );
  NOR2 U1037 ( .A(m1262), .B(m772), .OUT(N793) );
  INV U1038 ( .IN(\Samples[12][1] ), .OUT(m772) );
  NOR2 U1039 ( .A(m1262), .B(m773), .OUT(N792) );
  INV U1040 ( .IN(\Samples[12][0] ), .OUT(m773) );
  NOR2 U1041 ( .A(m1262), .B(m774), .OUT(N791) );
  INV U1042 ( .IN(\Samples[11][7] ), .OUT(m774) );
  NOR2 U1043 ( .A(m1262), .B(m775), .OUT(N790) );
  INV U1044 ( .IN(\Samples[11][6] ), .OUT(m775) );
  NOR2 U1045 ( .A(m1262), .B(m776), .OUT(N789) );
  INV U1046 ( .IN(\Samples[11][5] ), .OUT(m776) );
  NOR2 U1047 ( .A(m1262), .B(m777), .OUT(N788) );
  INV U1048 ( .IN(\Samples[11][4] ), .OUT(m777) );
  NOR2 U1049 ( .A(m1262), .B(m778), .OUT(N787) );
  INV U1050 ( .IN(\Samples[11][3] ), .OUT(m778) );
  NOR2 U1051 ( .A(m1262), .B(m779), .OUT(N786) );
  INV U1052 ( .IN(\Samples[11][2] ), .OUT(m779) );
  NOR2 U1053 ( .A(m1262), .B(m780), .OUT(N785) );
  INV U1054 ( .IN(\Samples[11][1] ), .OUT(m780) );
  NOR2 U1055 ( .A(m1262), .B(m781), .OUT(N784) );
  INV U1056 ( .IN(\Samples[11][0] ), .OUT(m781) );
  INV U1057 ( .IN(m782), .OUT(N920) );
  NAND2 U1058 ( .A(\Samples[10][7] ), .B(m1315), .OUT(m782) );
  INV U1059 ( .IN(m784), .OUT(N919) );
  NAND2 U1060 ( .A(\Samples[10][6] ), .B(m1315), .OUT(m784) );
  INV U1061 ( .IN(m785), .OUT(N918) );
  NAND2 U1062 ( .A(\Samples[10][5] ), .B(m1315), .OUT(m785) );
  INV U1063 ( .IN(m786), .OUT(N917) );
  NAND2 U1064 ( .A(\Samples[10][4] ), .B(m1314), .OUT(m786) );
  INV U1065 ( .IN(m787), .OUT(N916) );
  NAND2 U1066 ( .A(\Samples[10][3] ), .B(m1314), .OUT(m787) );
  INV U1067 ( .IN(m788), .OUT(N915) );
  NAND2 U1068 ( .A(\Samples[10][2] ), .B(m1314), .OUT(m788) );
  INV U1069 ( .IN(m789), .OUT(N914) );
  NAND2 U1070 ( .A(\Samples[10][1] ), .B(m1313), .OUT(m789) );
  INV U1071 ( .IN(m790), .OUT(N913) );
  NAND2 U1072 ( .A(\Samples[10][0] ), .B(m1313), .OUT(m790) );
  NOR2 U1073 ( .A(m1263), .B(m791), .OUT(N775) );
  INV U1074 ( .IN(\Samples[9][7] ), .OUT(m791) );
  NOR2 U1075 ( .A(m1263), .B(m792), .OUT(N774) );
  INV U1076 ( .IN(\Samples[9][6] ), .OUT(m792) );
  NOR2 U1077 ( .A(m1263), .B(m793), .OUT(N773) );
  INV U1078 ( .IN(\Samples[9][5] ), .OUT(m793) );
  NOR2 U1079 ( .A(m1263), .B(m794), .OUT(N772) );
  INV U1080 ( .IN(\Samples[9][4] ), .OUT(m794) );
  NOR2 U1081 ( .A(m1263), .B(m795), .OUT(N771) );
  INV U1082 ( .IN(\Samples[9][3] ), .OUT(m795) );
  NOR2 U1083 ( .A(m1263), .B(m796), .OUT(N770) );
  INV U1084 ( .IN(\Samples[9][2] ), .OUT(m796) );
  NOR2 U1085 ( .A(m1263), .B(m797), .OUT(N769) );
  INV U1086 ( .IN(\Samples[9][1] ), .OUT(m797) );
  NOR2 U1087 ( .A(m1263), .B(m798), .OUT(N768) );
  INV U1088 ( .IN(\Samples[9][0] ), .OUT(m798) );
  INV U1089 ( .IN(m799), .OUT(N901) );
  NAND2 U1090 ( .A(\Samples[8][7] ), .B(m1313), .OUT(m799) );
  INV U1091 ( .IN(m800), .OUT(N900) );
  NAND2 U1092 ( .A(\Samples[8][6] ), .B(m1312), .OUT(m800) );
  INV U1093 ( .IN(m801), .OUT(N899) );
  NAND2 U1094 ( .A(\Samples[8][5] ), .B(m1312), .OUT(m801) );
  INV U1095 ( .IN(m802), .OUT(N898) );
  NAND2 U1096 ( .A(\Samples[8][4] ), .B(m1312), .OUT(m802) );
  INV U1097 ( .IN(m803), .OUT(N897) );
  NAND2 U1098 ( .A(\Samples[8][3] ), .B(m1311), .OUT(m803) );
  INV U1099 ( .IN(m804), .OUT(N896) );
  NAND2 U1100 ( .A(\Samples[8][2] ), .B(m1311), .OUT(m804) );
  INV U1101 ( .IN(m805), .OUT(N895) );
  NAND2 U1102 ( .A(\Samples[8][1] ), .B(m1311), .OUT(m805) );
  INV U1103 ( .IN(m806), .OUT(N894) );
  NAND2 U1104 ( .A(\Samples[8][0] ), .B(m1310), .OUT(m806) );
  NOR2 U1105 ( .A(m1263), .B(m807), .OUT(N759) );
  INV U1106 ( .IN(\Samples[7][7] ), .OUT(m807) );
  NOR2 U1107 ( .A(m1263), .B(m808), .OUT(N758) );
  INV U1108 ( .IN(\Samples[7][6] ), .OUT(m808) );
  NOR2 U1109 ( .A(m1263), .B(m809), .OUT(N757) );
  INV U1110 ( .IN(\Samples[7][5] ), .OUT(m809) );
  NOR2 U1111 ( .A(m1263), .B(m810), .OUT(N756) );
  INV U1112 ( .IN(\Samples[7][4] ), .OUT(m810) );
  NOR2 U1113 ( .A(m1263), .B(m811), .OUT(N755) );
  INV U1114 ( .IN(\Samples[7][3] ), .OUT(m811) );
  NOR2 U1115 ( .A(m1264), .B(m812), .OUT(N754) );
  INV U1116 ( .IN(\Samples[7][2] ), .OUT(m812) );
  NOR2 U1117 ( .A(m1264), .B(m813), .OUT(N753) );
  INV U1118 ( .IN(\Samples[7][1] ), .OUT(m813) );
  NOR2 U1119 ( .A(m1264), .B(m814), .OUT(N752) );
  INV U1120 ( .IN(\Samples[7][0] ), .OUT(m814) );
  NOR2 U1121 ( .A(m1264), .B(m815), .OUT(N751) );
  INV U1122 ( .IN(\Samples[6][7] ), .OUT(m815) );
  NOR2 U1123 ( .A(m1264), .B(m816), .OUT(N750) );
  INV U1124 ( .IN(\Samples[6][6] ), .OUT(m816) );
  NOR2 U1125 ( .A(m1264), .B(m817), .OUT(N749) );
  INV U1126 ( .IN(\Samples[6][5] ), .OUT(m817) );
  NOR2 U1127 ( .A(m1264), .B(m818), .OUT(N748) );
  INV U1128 ( .IN(\Samples[6][4] ), .OUT(m818) );
  NOR2 U1129 ( .A(m1264), .B(m819), .OUT(N747) );
  INV U1130 ( .IN(\Samples[6][3] ), .OUT(m819) );
  NOR2 U1131 ( .A(m1264), .B(m820), .OUT(N746) );
  INV U1132 ( .IN(\Samples[6][2] ), .OUT(m820) );
  NOR2 U1133 ( .A(m1264), .B(m821), .OUT(N745) );
  INV U1134 ( .IN(\Samples[6][1] ), .OUT(m821) );
  NOR2 U1135 ( .A(m1264), .B(m822), .OUT(N744) );
  INV U1136 ( .IN(\Samples[6][0] ), .OUT(m822) );
  INV U1137 ( .IN(m823), .OUT(N869) );
  NAND2 U1138 ( .A(\Samples[5][7] ), .B(m1310), .OUT(m823) );
  INV U1139 ( .IN(m824), .OUT(N868) );
  NAND2 U1140 ( .A(\Samples[5][6] ), .B(m1310), .OUT(m824) );
  INV U1141 ( .IN(m825), .OUT(N867) );
  NAND2 U1142 ( .A(\Samples[5][5] ), .B(m1309), .OUT(m825) );
  INV U1143 ( .IN(m826), .OUT(N866) );
  NAND2 U1144 ( .A(\Samples[5][4] ), .B(m1309), .OUT(m826) );
  INV U1145 ( .IN(m827), .OUT(N865) );
  NAND2 U1146 ( .A(\Samples[5][3] ), .B(m1309), .OUT(m827) );
  INV U1147 ( .IN(m828), .OUT(N864) );
  NAND2 U1148 ( .A(\Samples[5][2] ), .B(m1308), .OUT(m828) );
  INV U1149 ( .IN(m829), .OUT(N863) );
  NAND2 U1150 ( .A(\Samples[5][1] ), .B(m1308), .OUT(m829) );
  INV U1151 ( .IN(m830), .OUT(N862) );
  NAND2 U1152 ( .A(\Samples[5][0] ), .B(m1308), .OUT(m830) );
  NOR2 U1153 ( .A(m1264), .B(m831), .OUT(N735) );
  INV U1154 ( .IN(\Samples[4][7] ), .OUT(m831) );
  NOR2 U1155 ( .A(m1264), .B(m832), .OUT(N734) );
  INV U1156 ( .IN(\Samples[4][6] ), .OUT(m832) );
  NOR2 U1157 ( .A(m1265), .B(m833), .OUT(N733) );
  INV U1158 ( .IN(\Samples[4][5] ), .OUT(m833) );
  NOR2 U1159 ( .A(m1265), .B(m834), .OUT(N732) );
  INV U1160 ( .IN(\Samples[4][4] ), .OUT(m834) );
  NOR2 U1161 ( .A(m1265), .B(m835), .OUT(N731) );
  INV U1162 ( .IN(\Samples[4][3] ), .OUT(m835) );
  NOR2 U1163 ( .A(m1265), .B(m836), .OUT(N730) );
  INV U1164 ( .IN(\Samples[4][2] ), .OUT(m836) );
  NOR2 U1165 ( .A(m1265), .B(m837), .OUT(N729) );
  INV U1166 ( .IN(\Samples[4][1] ), .OUT(m837) );
  NOR2 U1167 ( .A(m1265), .B(m838), .OUT(N728) );
  INV U1168 ( .IN(\Samples[4][0] ), .OUT(m838) );
  INV U1169 ( .IN(m839), .OUT(N850) );
  NAND2 U1170 ( .A(\Samples[3][7] ), .B(m1307), .OUT(m839) );
  INV U1171 ( .IN(m840), .OUT(N849) );
  NAND2 U1172 ( .A(\Samples[3][6] ), .B(m1307), .OUT(m840) );
  INV U1173 ( .IN(m841), .OUT(N848) );
  NAND2 U1174 ( .A(\Samples[3][5] ), .B(m1307), .OUT(m841) );
  INV U1175 ( .IN(m842), .OUT(N847) );
  NAND2 U1176 ( .A(\Samples[3][4] ), .B(m1306), .OUT(m842) );
  INV U1177 ( .IN(m843), .OUT(N846) );
  NAND2 U1178 ( .A(\Samples[3][3] ), .B(m1306), .OUT(m843) );
  INV U1179 ( .IN(m844), .OUT(N845) );
  NAND2 U1180 ( .A(\Samples[3][2] ), .B(m1306), .OUT(m844) );
  INV U1181 ( .IN(m845), .OUT(N844) );
  NAND2 U1182 ( .A(\Samples[3][1] ), .B(m1305), .OUT(m845) );
  INV U1183 ( .IN(m846), .OUT(N843) );
  NAND2 U1184 ( .A(\Samples[3][0] ), .B(m1305), .OUT(m846) );
  NOR2 U1185 ( .A(m1265), .B(m847), .OUT(N719) );
  INV U1186 ( .IN(\Samples[2][7] ), .OUT(m847) );
  NOR2 U1187 ( .A(m1265), .B(m848), .OUT(N718) );
  INV U1188 ( .IN(\Samples[2][6] ), .OUT(m848) );
  NOR2 U1189 ( .A(m1265), .B(m849), .OUT(N717) );
  INV U1190 ( .IN(\Samples[2][5] ), .OUT(m849) );
  NOR2 U1191 ( .A(m1265), .B(m850), .OUT(N716) );
  INV U1192 ( .IN(\Samples[2][4] ), .OUT(m850) );
  NOR2 U1193 ( .A(m1265), .B(m851), .OUT(N715) );
  INV U1194 ( .IN(\Samples[2][3] ), .OUT(m851) );
  NOR2 U1195 ( .A(m1265), .B(m852), .OUT(N714) );
  INV U1196 ( .IN(\Samples[2][2] ), .OUT(m852) );
  NOR2 U1197 ( .A(m1265), .B(m853), .OUT(N713) );
  INV U1198 ( .IN(\Samples[2][1] ), .OUT(m853) );
  NOR2 U1199 ( .A(m1266), .B(m854), .OUT(N712) );
  INV U1200 ( .IN(\Samples[2][0] ), .OUT(m854) );
  NOR2 U1201 ( .A(m1266), .B(m855), .OUT(N711) );
  INV U1202 ( .IN(\Samples[1][7] ), .OUT(m855) );
  NOR2 U1203 ( .A(m1266), .B(m856), .OUT(N710) );
  INV U1204 ( .IN(\Samples[1][6] ), .OUT(m856) );
  NOR2 U1205 ( .A(m1266), .B(m857), .OUT(N709) );
  INV U1206 ( .IN(\Samples[1][5] ), .OUT(m857) );
  NOR2 U1207 ( .A(m1266), .B(m858), .OUT(N708) );
  INV U1208 ( .IN(\Samples[1][4] ), .OUT(m858) );
  NOR2 U1209 ( .A(m1266), .B(m859), .OUT(N707) );
  INV U1210 ( .IN(\Samples[1][3] ), .OUT(m859) );
  NOR2 U1211 ( .A(m1266), .B(m860), .OUT(N706) );
  INV U1212 ( .IN(\Samples[1][2] ), .OUT(m860) );
  NOR2 U1213 ( .A(m1266), .B(m861), .OUT(N705) );
  INV U1214 ( .IN(\Samples[1][1] ), .OUT(m861) );
  NOR2 U1215 ( .A(m1266), .B(m862), .OUT(N704) );
  INV U1216 ( .IN(\Samples[1][0] ), .OUT(m862) );
  INV U1217 ( .IN(m863), .OUT(N818) );
  NAND2 U1218 ( .A(\Samples[0][7] ), .B(m1305), .OUT(m863) );
  INV U1219 ( .IN(m864), .OUT(N817) );
  NAND2 U1220 ( .A(\Samples[0][6] ), .B(m1304), .OUT(m864) );
  INV U1221 ( .IN(m865), .OUT(N816) );
  NAND2 U1222 ( .A(\Samples[0][5] ), .B(m1304), .OUT(m865) );
  INV U1223 ( .IN(m866), .OUT(N815) );
  NAND2 U1224 ( .A(\Samples[0][4] ), .B(m1304), .OUT(m866) );
  INV U1225 ( .IN(m867), .OUT(N814) );
  NAND2 U1226 ( .A(\Samples[0][3] ), .B(m1303), .OUT(m867) );
  INV U1227 ( .IN(m868), .OUT(N813) );
  NAND2 U1228 ( .A(\Samples[0][2] ), .B(m1303), .OUT(m868) );
  INV U1229 ( .IN(m869), .OUT(N812) );
  NAND2 U1230 ( .A(\Samples[0][1] ), .B(m1303), .OUT(m869) );
  INV U1231 ( .IN(m870), .OUT(N811) );
  NAND2 U1232 ( .A(\Samples[0][0] ), .B(m1302), .OUT(m870) );
  NOR2 U1234 ( .A(m1266), .B(m871), .OUT(N695) );
  INV U1235 ( .IN(Data_in[7]), .OUT(m871) );
  NOR2 U1236 ( .A(m1266), .B(m872), .OUT(N694) );
  INV U1237 ( .IN(Data_in[6]), .OUT(m872) );
  NOR2 U1238 ( .A(m1266), .B(m873), .OUT(N693) );
  INV U1239 ( .IN(Data_in[5]), .OUT(m873) );
  NOR2 U1240 ( .A(m1266), .B(m874), .OUT(N692) );
  INV U1241 ( .IN(Data_in[4]), .OUT(m874) );
  NOR2 U1242 ( .A(m1267), .B(m875), .OUT(N691) );
  INV U1243 ( .IN(Data_in[3]), .OUT(m875) );
  NOR2 U1244 ( .A(m1267), .B(m876), .OUT(N690) );
  INV U1245 ( .IN(Data_in[2]), .OUT(m876) );
  NOR2 U1246 ( .A(m1267), .B(m877), .OUT(N689) );
  INV U1247 ( .IN(Data_in[1]), .OUT(m877) );
  NOR2 U1248 ( .A(m1267), .B(m878), .OUT(N688) );
  INV U1249 ( .IN(Data_in[0]), .OUT(m878) );
  NOR2 U1250 ( .A(m1267), .B(m879), .OUT(N687) );
  INV U1251 ( .IN(N387), .OUT(m879) );
  NOR2 U1252 ( .A(m1267), .B(m880), .OUT(N686) );
  INV U1253 ( .IN(N386), .OUT(m880) );
  NOR2 U1254 ( .A(m1267), .B(m881), .OUT(N685) );
  INV U1255 ( .IN(N385), .OUT(m881) );
  NOR2 U1256 ( .A(m1267), .B(m882), .OUT(N684) );
  INV U1257 ( .IN(N384), .OUT(m882) );
  NOR2 U1258 ( .A(m1267), .B(m883), .OUT(N683) );
  INV U1259 ( .IN(N383), .OUT(m883) );
  NOR2 U1260 ( .A(m1267), .B(m884), .OUT(N682) );
  INV U1261 ( .IN(N382), .OUT(m884) );
  NOR2 U1262 ( .A(m1267), .B(m885), .OUT(N681) );
  INV U1263 ( .IN(N381), .OUT(m885) );
  NOR2 U1264 ( .A(m1267), .B(m886), .OUT(N680) );
  INV U1265 ( .IN(N380), .OUT(m886) );
  NOR2 U1266 ( .A(m1267), .B(m887), .OUT(N679) );
  INV U1267 ( .IN(N379), .OUT(m887) );
  NOR2 U1268 ( .A(m1268), .B(m888), .OUT(N678) );
  INV U1269 ( .IN(N378), .OUT(m888) );
  NOR2 U1270 ( .A(m1268), .B(m889), .OUT(N677) );
  INV U1271 ( .IN(N377), .OUT(m889) );
  NOR2 U1272 ( .A(m1268), .B(m890), .OUT(N676) );
  INV U1273 ( .IN(N376), .OUT(m890) );
  NOR2 U1274 ( .A(m1268), .B(m891), .OUT(N675) );
  INV U1275 ( .IN(N375), .OUT(m891) );
  NOR2 U1276 ( .A(m1268), .B(m892), .OUT(N674) );
  INV U1277 ( .IN(N374), .OUT(m892) );
  NOR2 U1278 ( .A(m1268), .B(m893), .OUT(N673) );
  INV U1279 ( .IN(N373), .OUT(m893) );
  NOR2 U1280 ( .A(m1268), .B(m894), .OUT(N672) );
  INV U1281 ( .IN(N372), .OUT(m894) );
  NOR2 U1282 ( .A(m1268), .B(m895), .OUT(N671) );
  INV U1283 ( .IN(N371), .OUT(m895) );
  NOR2 U1284 ( .A(m1268), .B(m896), .OUT(N670) );
  INV U1285 ( .IN(N370), .OUT(m896) );
  NOR2 U1286 ( .A(m1268), .B(m897), .OUT(N669) );
  INV U1287 ( .IN(N369), .OUT(m897) );
  NOR2 U1288 ( .A(m1268), .B(m898), .OUT(N668) );
  INV U1289 ( .IN(N368), .OUT(m898) );
  NOR2 U1290 ( .A(m1268), .B(m899), .OUT(N667) );
  INV U1291 ( .IN(N367), .OUT(m899) );
  NOR2 U1292 ( .A(m1268), .B(m900), .OUT(N666) );
  INV U1293 ( .IN(N366), .OUT(m900) );
  NOR2 U1294 ( .A(m1269), .B(m901), .OUT(N665) );
  INV U1295 ( .IN(N365), .OUT(m901) );
  NOR2 U1296 ( .A(m1269), .B(m902), .OUT(N664) );
  INV U1297 ( .IN(N364), .OUT(m902) );
  NOR2 U1298 ( .A(m1269), .B(m903), .OUT(N663) );
  INV U1299 ( .IN(N363), .OUT(m903) );
  NOR2 U1300 ( .A(m1269), .B(m904), .OUT(N662) );
  INV U1301 ( .IN(N362), .OUT(m904) );
  NOR2 U1302 ( .A(m1269), .B(m905), .OUT(N661) );
  INV U1303 ( .IN(N361), .OUT(m905) );
  NOR2 U1304 ( .A(m1269), .B(m906), .OUT(N660) );
  INV U1305 ( .IN(N360), .OUT(m906) );
  NOR2 U1306 ( .A(m1269), .B(m907), .OUT(N659) );
  INV U1307 ( .IN(N359), .OUT(m907) );
  NOR2 U1308 ( .A(m1269), .B(m908), .OUT(N658) );
  INV U1309 ( .IN(N358), .OUT(m908) );
  NOR2 U1310 ( .A(m1269), .B(m909), .OUT(N657) );
  INV U1311 ( .IN(N357), .OUT(m909) );
  NOR2 U1312 ( .A(m1269), .B(m910), .OUT(N656) );
  INV U1313 ( .IN(N356), .OUT(m910) );
  NOR2 U1314 ( .A(m1269), .B(m911), .OUT(N655) );
  INV U1315 ( .IN(N355), .OUT(m911) );
  NOR2 U1316 ( .A(m1269), .B(m912), .OUT(N654) );
  INV U1317 ( .IN(N354), .OUT(m912) );
  NOR2 U1318 ( .A(m1269), .B(m913), .OUT(N653) );
  INV U1319 ( .IN(N353), .OUT(m913) );
  NOR2 U1320 ( .A(m1270), .B(m914), .OUT(N652) );
  INV U1321 ( .IN(N352), .OUT(m914) );
  NOR2 U1322 ( .A(m1270), .B(m915), .OUT(N651) );
  INV U1323 ( .IN(N351), .OUT(m915) );
  NOR2 U1324 ( .A(m1270), .B(m916), .OUT(N650) );
  INV U1325 ( .IN(N350), .OUT(m916) );
  NOR2 U1326 ( .A(m1270), .B(m917), .OUT(N649) );
  INV U1327 ( .IN(N349), .OUT(m917) );
  NOR2 U1328 ( .A(m1270), .B(m918), .OUT(N648) );
  INV U1329 ( .IN(N348), .OUT(m918) );
  NOR2 U1330 ( .A(m1270), .B(m919), .OUT(N647) );
  INV U1331 ( .IN(N347), .OUT(m919) );
  NOR2 U1332 ( .A(m1270), .B(m920), .OUT(N646) );
  INV U1333 ( .IN(N346), .OUT(m920) );
  NOR2 U1334 ( .A(m1270), .B(m921), .OUT(N645) );
  INV U1335 ( .IN(N345), .OUT(m921) );
  NOR2 U1336 ( .A(m1270), .B(m922), .OUT(N644) );
  INV U1337 ( .IN(N344), .OUT(m922) );
  NOR2 U1338 ( .A(m1270), .B(m923), .OUT(N643) );
  INV U1339 ( .IN(N343), .OUT(m923) );
  NOR2 U1340 ( .A(m1270), .B(m924), .OUT(N642) );
  INV U1341 ( .IN(N342), .OUT(m924) );
  NOR2 U1342 ( .A(m1270), .B(m925), .OUT(N641) );
  INV U1343 ( .IN(N341), .OUT(m925) );
  NOR2 U1344 ( .A(m1270), .B(m926), .OUT(N640) );
  INV U1345 ( .IN(N340), .OUT(m926) );
  NOR2 U1346 ( .A(m1271), .B(m927), .OUT(N639) );
  INV U1347 ( .IN(N339), .OUT(m927) );
  NOR2 U1348 ( .A(m1271), .B(m928), .OUT(N638) );
  INV U1349 ( .IN(N338), .OUT(m928) );
  NOR2 U1350 ( .A(m1271), .B(m929), .OUT(N637) );
  INV U1351 ( .IN(N337), .OUT(m929) );
  NOR2 U1352 ( .A(m1271), .B(m930), .OUT(N636) );
  INV U1353 ( .IN(N336), .OUT(m930) );
  NOR2 U1354 ( .A(m1271), .B(m931), .OUT(N635) );
  INV U1355 ( .IN(N335), .OUT(m931) );
  NOR2 U1356 ( .A(m1271), .B(m932), .OUT(N634) );
  INV U1357 ( .IN(N334), .OUT(m932) );
  NOR2 U1358 ( .A(m1271), .B(m933), .OUT(N633) );
  INV U1359 ( .IN(N333), .OUT(m933) );
  NOR2 U1360 ( .A(m1271), .B(m934), .OUT(N632) );
  INV U1361 ( .IN(N332), .OUT(m934) );
  NOR2 U1362 ( .A(m1271), .B(m935), .OUT(N631) );
  INV U1363 ( .IN(N331), .OUT(m935) );
  NOR2 U1364 ( .A(m1271), .B(m936), .OUT(N630) );
  INV U1365 ( .IN(N330), .OUT(m936) );
  NOR2 U1366 ( .A(m1271), .B(m937), .OUT(N629) );
  INV U1367 ( .IN(N329), .OUT(m937) );
  NOR2 U1368 ( .A(m1271), .B(m938), .OUT(N628) );
  INV U1369 ( .IN(N328), .OUT(m938) );
  NOR2 U1370 ( .A(m1271), .B(m939), .OUT(N627) );
  INV U1371 ( .IN(N327), .OUT(m939) );
  NOR2 U1372 ( .A(m1272), .B(m940), .OUT(N626) );
  INV U1373 ( .IN(N326), .OUT(m940) );
  NOR2 U1374 ( .A(m1272), .B(m941), .OUT(N625) );
  INV U1375 ( .IN(N325), .OUT(m941) );
  NOR2 U1376 ( .A(m1272), .B(m942), .OUT(N624) );
  INV U1377 ( .IN(N324), .OUT(m942) );
  NOR2 U1378 ( .A(m1272), .B(m943), .OUT(N623) );
  INV U1379 ( .IN(N323), .OUT(m943) );
  NOR2 U1380 ( .A(m1272), .B(m944), .OUT(N622) );
  INV U1381 ( .IN(N322), .OUT(m944) );
  NOR2 U1382 ( .A(m1272), .B(m945), .OUT(N621) );
  INV U1383 ( .IN(N321), .OUT(m945) );
  NOR2 U1384 ( .A(m1272), .B(m946), .OUT(N620) );
  INV U1385 ( .IN(N320), .OUT(m946) );
  NOR2 U1386 ( .A(m1272), .B(m947), .OUT(N619) );
  INV U1387 ( .IN(N319), .OUT(m947) );
  NOR2 U1388 ( .A(m1272), .B(m948), .OUT(N618) );
  INV U1389 ( .IN(N318), .OUT(m948) );
  NOR2 U1390 ( .A(m1272), .B(m949), .OUT(N617) );
  INV U1391 ( .IN(N317), .OUT(m949) );
  NOR2 U1392 ( .A(m1272), .B(m950), .OUT(N616) );
  INV U1393 ( .IN(N316), .OUT(m950) );
  NOR2 U1394 ( .A(m1272), .B(m951), .OUT(N615) );
  INV U1395 ( .IN(N315), .OUT(m951) );
  NOR2 U1396 ( .A(m1272), .B(m952), .OUT(N614) );
  INV U1397 ( .IN(N314), .OUT(m952) );
  NOR2 U1398 ( .A(m1273), .B(m953), .OUT(N613) );
  INV U1399 ( .IN(N313), .OUT(m953) );
  NOR2 U1400 ( .A(m1273), .B(m954), .OUT(N612) );
  INV U1401 ( .IN(N312), .OUT(m954) );
  NOR2 U1402 ( .A(m1273), .B(m955), .OUT(N611) );
  INV U1403 ( .IN(N311), .OUT(m955) );
  NOR2 U1404 ( .A(m1273), .B(m956), .OUT(N610) );
  INV U1405 ( .IN(N310), .OUT(m956) );
  NOR2 U1406 ( .A(m1273), .B(m957), .OUT(N609) );
  INV U1407 ( .IN(N309), .OUT(m957) );
  NOR2 U1408 ( .A(m1273), .B(m958), .OUT(N608) );
  INV U1409 ( .IN(N308), .OUT(m958) );
  NOR2 U1410 ( .A(m1273), .B(m959), .OUT(N607) );
  INV U1411 ( .IN(N307), .OUT(m959) );
  NOR2 U1412 ( .A(m1273), .B(m960), .OUT(N606) );
  INV U1413 ( .IN(N306), .OUT(m960) );
  NOR2 U1414 ( .A(m1273), .B(m961), .OUT(N605) );
  INV U1415 ( .IN(N305), .OUT(m961) );
  NOR2 U1416 ( .A(m1273), .B(m962), .OUT(N604) );
  INV U1417 ( .IN(N304), .OUT(m962) );
  NOR2 U1418 ( .A(m1273), .B(m963), .OUT(N603) );
  INV U1419 ( .IN(N303), .OUT(m963) );
  NOR2 U1420 ( .A(m1273), .B(m964), .OUT(N602) );
  INV U1421 ( .IN(N302), .OUT(m964) );
  NOR2 U1422 ( .A(m1273), .B(m965), .OUT(N601) );
  INV U1423 ( .IN(N301), .OUT(m965) );
  NOR2 U1424 ( .A(m1274), .B(m966), .OUT(N600) );
  INV U1425 ( .IN(N300), .OUT(m966) );
  NOR2 U1426 ( .A(m1274), .B(m967), .OUT(N599) );
  INV U1427 ( .IN(N299), .OUT(m967) );
  NOR2 U1428 ( .A(m1274), .B(m968), .OUT(N598) );
  INV U1429 ( .IN(N298), .OUT(m968) );
  NOR2 U1430 ( .A(m1274), .B(m969), .OUT(N597) );
  INV U1431 ( .IN(N297), .OUT(m969) );
  NOR2 U1432 ( .A(m1274), .B(m970), .OUT(N596) );
  INV U1433 ( .IN(N296), .OUT(m970) );
  NOR2 U1434 ( .A(m1274), .B(m971), .OUT(N595) );
  INV U1435 ( .IN(N295), .OUT(m971) );
  NOR2 U1436 ( .A(m1274), .B(m972), .OUT(N594) );
  INV U1437 ( .IN(N294), .OUT(m972) );
  NOR2 U1438 ( .A(m1274), .B(m973), .OUT(N593) );
  INV U1439 ( .IN(N293), .OUT(m973) );
  NOR2 U1440 ( .A(m1274), .B(m974), .OUT(N592) );
  INV U1441 ( .IN(N292), .OUT(m974) );
  NOR2 U1442 ( .A(m1274), .B(m975), .OUT(N591) );
  INV U1443 ( .IN(N291), .OUT(m975) );
  NOR2 U1444 ( .A(m1274), .B(m976), .OUT(N590) );
  INV U1445 ( .IN(N290), .OUT(m976) );
  NOR2 U1446 ( .A(m1274), .B(m977), .OUT(N589) );
  INV U1447 ( .IN(N289), .OUT(m977) );
  NOR2 U1448 ( .A(m1274), .B(m978), .OUT(N588) );
  INV U1449 ( .IN(N288), .OUT(m978) );
  NOR2 U1450 ( .A(m1275), .B(m979), .OUT(N587) );
  INV U1451 ( .IN(N287), .OUT(m979) );
  NOR2 U1452 ( .A(m1275), .B(m980), .OUT(N586) );
  INV U1453 ( .IN(N286), .OUT(m980) );
  NOR2 U1454 ( .A(m1275), .B(m981), .OUT(N585) );
  INV U1455 ( .IN(N285), .OUT(m981) );
  NOR2 U1456 ( .A(m1275), .B(m982), .OUT(N584) );
  INV U1457 ( .IN(N284), .OUT(m982) );
  NOR2 U1458 ( .A(m1275), .B(m983), .OUT(N583) );
  INV U1459 ( .IN(N283), .OUT(m983) );
  NOR2 U1460 ( .A(m1275), .B(m984), .OUT(N582) );
  INV U1461 ( .IN(N282), .OUT(m984) );
  NOR2 U1462 ( .A(m1275), .B(m985), .OUT(N581) );
  INV U1463 ( .IN(N281), .OUT(m985) );
  NOR2 U1464 ( .A(m1275), .B(m986), .OUT(N580) );
  INV U1465 ( .IN(N280), .OUT(m986) );
  NOR2 U1466 ( .A(m1275), .B(m987), .OUT(N579) );
  INV U1467 ( .IN(N279), .OUT(m987) );
  NOR2 U1468 ( .A(m1275), .B(m988), .OUT(N578) );
  INV U1469 ( .IN(N278), .OUT(m988) );
  NOR2 U1470 ( .A(m1275), .B(m989), .OUT(N577) );
  INV U1471 ( .IN(N277), .OUT(m989) );
  NOR2 U1472 ( .A(m1275), .B(m990), .OUT(N576) );
  INV U1473 ( .IN(N276), .OUT(m990) );
  NOR2 U1474 ( .A(m1275), .B(m991), .OUT(N575) );
  INV U1475 ( .IN(N275), .OUT(m991) );
  NOR2 U1476 ( .A(m1276), .B(m992), .OUT(N574) );
  INV U1477 ( .IN(N274), .OUT(m992) );
  NOR2 U1478 ( .A(m1276), .B(m993), .OUT(N573) );
  INV U1479 ( .IN(N273), .OUT(m993) );
  NOR2 U1480 ( .A(m1276), .B(m994), .OUT(N572) );
  INV U1481 ( .IN(N272), .OUT(m994) );
  NOR2 U1482 ( .A(m1276), .B(m995), .OUT(N571) );
  INV U1483 ( .IN(N271), .OUT(m995) );
  NOR2 U1484 ( .A(m1276), .B(m996), .OUT(N570) );
  INV U1485 ( .IN(N270), .OUT(m996) );
  NOR2 U1486 ( .A(m1276), .B(m997), .OUT(N569) );
  INV U1487 ( .IN(N269), .OUT(m997) );
  NOR2 U1488 ( .A(m1276), .B(m998), .OUT(N568) );
  INV U1489 ( .IN(N268), .OUT(m998) );
  NOR2 U1490 ( .A(m1276), .B(m999), .OUT(N567) );
  INV U1491 ( .IN(N267), .OUT(m999) );
  NOR2 U1492 ( .A(m1276), .B(m1000), .OUT(N566) );
  INV U1493 ( .IN(N266), .OUT(m1000) );
  NOR2 U1494 ( .A(m1276), .B(m1001), .OUT(N565) );
  INV U1495 ( .IN(N265), .OUT(m1001) );
  NOR2 U1496 ( .A(m1276), .B(m1002), .OUT(N564) );
  INV U1497 ( .IN(N264), .OUT(m1002) );
  NOR2 U1498 ( .A(m1276), .B(m1003), .OUT(N563) );
  INV U1499 ( .IN(N263), .OUT(m1003) );
  NOR2 U1500 ( .A(m1276), .B(m1004), .OUT(N562) );
  INV U1501 ( .IN(N262), .OUT(m1004) );
  NOR2 U1502 ( .A(m1277), .B(m1005), .OUT(N561) );
  INV U1503 ( .IN(N261), .OUT(m1005) );
  NOR2 U1504 ( .A(m1277), .B(m1006), .OUT(N560) );
  INV U1505 ( .IN(N260), .OUT(m1006) );
  NOR2 U1506 ( .A(m1277), .B(m1007), .OUT(N559) );
  INV U1507 ( .IN(N259), .OUT(m1007) );
  NOR2 U1508 ( .A(m1277), .B(m1008), .OUT(N558) );
  INV U1509 ( .IN(N258), .OUT(m1008) );
  NOR2 U1510 ( .A(m1277), .B(m1009), .OUT(N557) );
  INV U1511 ( .IN(N257), .OUT(m1009) );
  NOR2 U1512 ( .A(m1277), .B(m1010), .OUT(N556) );
  INV U1513 ( .IN(N256), .OUT(m1010) );
  NOR2 U1514 ( .A(m1277), .B(m1011), .OUT(N555) );
  INV U1515 ( .IN(N255), .OUT(m1011) );
  NOR2 U1516 ( .A(m1277), .B(m1012), .OUT(N554) );
  INV U1517 ( .IN(N254), .OUT(m1012) );
  NOR2 U1518 ( .A(m1277), .B(m1013), .OUT(N553) );
  INV U1519 ( .IN(N253), .OUT(m1013) );
  NOR2 U1520 ( .A(m1277), .B(m1014), .OUT(N552) );
  INV U1521 ( .IN(N252), .OUT(m1014) );
  NOR2 U1522 ( .A(m1277), .B(m1015), .OUT(N551) );
  INV U1523 ( .IN(N251), .OUT(m1015) );
  NOR2 U1524 ( .A(m1277), .B(m1016), .OUT(N550) );
  INV U1525 ( .IN(N250), .OUT(m1016) );
  NOR2 U1526 ( .A(m1277), .B(m1017), .OUT(N549) );
  INV U1527 ( .IN(N249), .OUT(m1017) );
  NOR2 U1528 ( .A(m1278), .B(m1018), .OUT(N548) );
  INV U1529 ( .IN(N248), .OUT(m1018) );
  NOR2 U1530 ( .A(m1278), .B(m1019), .OUT(N547) );
  INV U1531 ( .IN(N247), .OUT(m1019) );
  NOR2 U1532 ( .A(m1278), .B(m1020), .OUT(N546) );
  INV U1533 ( .IN(N246), .OUT(m1020) );
  NOR2 U1534 ( .A(m1278), .B(m1021), .OUT(N545) );
  INV U1535 ( .IN(N245), .OUT(m1021) );
  NOR2 U1536 ( .A(m1278), .B(m1022), .OUT(N544) );
  INV U1537 ( .IN(N244), .OUT(m1022) );
  NOR2 U1538 ( .A(m1278), .B(m1023), .OUT(N543) );
  INV U1539 ( .IN(N243), .OUT(m1023) );
  NOR2 U1540 ( .A(m1278), .B(m1024), .OUT(N542) );
  INV U1541 ( .IN(N242), .OUT(m1024) );
  NOR2 U1542 ( .A(m1278), .B(m1025), .OUT(N541) );
  INV U1543 ( .IN(N241), .OUT(m1025) );
  NOR2 U1544 ( .A(m1278), .B(m1026), .OUT(N540) );
  INV U1545 ( .IN(N240), .OUT(m1026) );
  NOR2 U1546 ( .A(m1278), .B(m1027), .OUT(N539) );
  INV U1547 ( .IN(N239), .OUT(m1027) );
  NOR2 U1548 ( .A(m1278), .B(m1028), .OUT(N538) );
  INV U1549 ( .IN(N238), .OUT(m1028) );
  NOR2 U1550 ( .A(m1278), .B(m1029), .OUT(N537) );
  INV U1551 ( .IN(N237), .OUT(m1029) );
  NOR2 U1552 ( .A(m1278), .B(m1030), .OUT(N536) );
  INV U1553 ( .IN(N236), .OUT(m1030) );
  NOR2 U1554 ( .A(m1279), .B(m1031), .OUT(N535) );
  INV U1555 ( .IN(N235), .OUT(m1031) );
  NOR2 U1556 ( .A(m1279), .B(m1032), .OUT(N534) );
  INV U1557 ( .IN(N234), .OUT(m1032) );
  NOR2 U1558 ( .A(m1279), .B(m1033), .OUT(N533) );
  INV U1559 ( .IN(N233), .OUT(m1033) );
  NOR2 U1560 ( .A(m1279), .B(m1034), .OUT(N532) );
  INV U1561 ( .IN(N232), .OUT(m1034) );
  NOR2 U1562 ( .A(m1279), .B(m1035), .OUT(N531) );
  INV U1563 ( .IN(N231), .OUT(m1035) );
  NOR2 U1564 ( .A(m1279), .B(m1036), .OUT(N530) );
  INV U1565 ( .IN(N230), .OUT(m1036) );
  NOR2 U1566 ( .A(m1279), .B(m1037), .OUT(N529) );
  INV U1567 ( .IN(N229), .OUT(m1037) );
  NOR2 U1568 ( .A(m1279), .B(m1038), .OUT(N528) );
  INV U1569 ( .IN(N228), .OUT(m1038) );
  NOR2 U1570 ( .A(m1279), .B(m1039), .OUT(N527) );
  INV U1571 ( .IN(N227), .OUT(m1039) );
  NOR2 U1572 ( .A(m1279), .B(m1040), .OUT(N526) );
  INV U1573 ( .IN(N226), .OUT(m1040) );
  NOR2 U1574 ( .A(m1279), .B(m1041), .OUT(N525) );
  INV U1575 ( .IN(N225), .OUT(m1041) );
  NOR2 U1576 ( .A(m1279), .B(m1042), .OUT(N524) );
  INV U1577 ( .IN(N224), .OUT(m1042) );
  NOR2 U1578 ( .A(m1279), .B(m1043), .OUT(N523) );
  INV U1579 ( .IN(N223), .OUT(m1043) );
  NOR2 U1580 ( .A(m1280), .B(m1044), .OUT(N522) );
  INV U1581 ( .IN(N222), .OUT(m1044) );
  NOR2 U1582 ( .A(m1280), .B(m1045), .OUT(N521) );
  INV U1583 ( .IN(N221), .OUT(m1045) );
  NOR2 U1584 ( .A(m1280), .B(m1046), .OUT(N520) );
  INV U1585 ( .IN(N220), .OUT(m1046) );
  NOR2 U1586 ( .A(m1280), .B(m1047), .OUT(N519) );
  INV U1587 ( .IN(N219), .OUT(m1047) );
  NOR2 U1588 ( .A(m1280), .B(m1048), .OUT(N518) );
  INV U1589 ( .IN(N218), .OUT(m1048) );
  NOR2 U1590 ( .A(m1280), .B(m1049), .OUT(N517) );
  INV U1591 ( .IN(N217), .OUT(m1049) );
  NOR2 U1592 ( .A(m1280), .B(m1050), .OUT(N516) );
  INV U1593 ( .IN(N216), .OUT(m1050) );
  NOR2 U1594 ( .A(m1280), .B(m1051), .OUT(N515) );
  INV U1595 ( .IN(N215), .OUT(m1051) );
  NOR2 U1596 ( .A(m1280), .B(m1052), .OUT(N514) );
  INV U1597 ( .IN(N214), .OUT(m1052) );
  NOR2 U1598 ( .A(m1280), .B(m1053), .OUT(N513) );
  INV U1599 ( .IN(N213), .OUT(m1053) );
  NOR2 U1600 ( .A(m1280), .B(m1054), .OUT(N512) );
  INV U1601 ( .IN(N212), .OUT(m1054) );
  NOR2 U1602 ( .A(m1280), .B(m1055), .OUT(N511) );
  INV U1603 ( .IN(N211), .OUT(m1055) );
  NOR2 U1604 ( .A(m1280), .B(m1056), .OUT(N510) );
  INV U1605 ( .IN(N210), .OUT(m1056) );
  NOR2 U1606 ( .A(m1281), .B(m1057), .OUT(N509) );
  INV U1607 ( .IN(N209), .OUT(m1057) );
  NOR2 U1608 ( .A(m1281), .B(m1058), .OUT(N508) );
  INV U1609 ( .IN(N208), .OUT(m1058) );
  NOR2 U1610 ( .A(m1281), .B(m1059), .OUT(N507) );
  INV U1611 ( .IN(N207), .OUT(m1059) );
  NOR2 U1612 ( .A(m1281), .B(m1060), .OUT(N506) );
  INV U1613 ( .IN(N206), .OUT(m1060) );
  NOR2 U1614 ( .A(m1281), .B(m1061), .OUT(N505) );
  INV U1615 ( .IN(N205), .OUT(m1061) );
  NOR2 U1616 ( .A(m1281), .B(m1062), .OUT(N504) );
  INV U1617 ( .IN(N204), .OUT(m1062) );
  NOR2 U1618 ( .A(m1281), .B(m1063), .OUT(N503) );
  INV U1619 ( .IN(N203), .OUT(m1063) );
  NOR2 U1620 ( .A(m1281), .B(m1064), .OUT(N502) );
  INV U1621 ( .IN(N202), .OUT(m1064) );
  NOR2 U1622 ( .A(m1281), .B(m1065), .OUT(N501) );
  INV U1623 ( .IN(N201), .OUT(m1065) );
  NOR2 U1624 ( .A(m1281), .B(m1066), .OUT(N500) );
  INV U1625 ( .IN(N200), .OUT(m1066) );
  NOR2 U1626 ( .A(m1281), .B(m1067), .OUT(N499) );
  INV U1627 ( .IN(N199), .OUT(m1067) );
  NOR2 U1628 ( .A(m1281), .B(m1068), .OUT(N498) );
  INV U1629 ( .IN(N198), .OUT(m1068) );
  NOR2 U1630 ( .A(m1281), .B(m1069), .OUT(N497) );
  INV U1631 ( .IN(N197), .OUT(m1069) );
  NOR2 U1632 ( .A(m1282), .B(m1070), .OUT(N496) );
  INV U1633 ( .IN(N196), .OUT(m1070) );
  NOR2 U1634 ( .A(m1282), .B(m1071), .OUT(N495) );
  INV U1635 ( .IN(N195), .OUT(m1071) );
  NOR2 U1636 ( .A(m1282), .B(m1072), .OUT(N494) );
  INV U1637 ( .IN(N194), .OUT(m1072) );
  NOR2 U1638 ( .A(m1282), .B(m1073), .OUT(N493) );
  INV U1639 ( .IN(N193), .OUT(m1073) );
  NOR2 U1640 ( .A(m1282), .B(m1074), .OUT(N492) );
  INV U1641 ( .IN(N192), .OUT(m1074) );
  NOR2 U1642 ( .A(m1282), .B(m1075), .OUT(N491) );
  INV U1643 ( .IN(N191), .OUT(m1075) );
  NOR2 U1644 ( .A(m1282), .B(m1076), .OUT(N490) );
  INV U1645 ( .IN(N190), .OUT(m1076) );
  NOR2 U1646 ( .A(m1282), .B(m1077), .OUT(N489) );
  INV U1647 ( .IN(N189), .OUT(m1077) );
  NOR2 U1648 ( .A(m1282), .B(m1078), .OUT(N488) );
  INV U1649 ( .IN(N188), .OUT(m1078) );
  NOR2 U1650 ( .A(m1282), .B(m1079), .OUT(N487) );
  INV U1651 ( .IN(N187), .OUT(m1079) );
  NOR2 U1652 ( .A(m1282), .B(m1080), .OUT(N486) );
  INV U1653 ( .IN(N186), .OUT(m1080) );
  NOR2 U1654 ( .A(m1282), .B(m1081), .OUT(N485) );
  INV U1655 ( .IN(N185), .OUT(m1081) );
  NOR2 U1656 ( .A(m1282), .B(m1082), .OUT(N484) );
  INV U1657 ( .IN(N184), .OUT(m1082) );
  NOR2 U1658 ( .A(m1283), .B(m1083), .OUT(N483) );
  INV U1659 ( .IN(N183), .OUT(m1083) );
  NOR2 U1660 ( .A(m1283), .B(m1084), .OUT(N482) );
  INV U1661 ( .IN(N182), .OUT(m1084) );
  NOR2 U1662 ( .A(m1283), .B(m1085), .OUT(N481) );
  INV U1663 ( .IN(N181), .OUT(m1085) );
  NOR2 U1664 ( .A(m1283), .B(m1086), .OUT(N480) );
  INV U1665 ( .IN(N180), .OUT(m1086) );
  NOR2 U1666 ( .A(m1283), .B(m1087), .OUT(N479) );
  INV U1667 ( .IN(N179), .OUT(m1087) );
  NOR2 U1668 ( .A(m1283), .B(m1088), .OUT(N478) );
  INV U1669 ( .IN(N178), .OUT(m1088) );
  NOR2 U1670 ( .A(m1283), .B(m1089), .OUT(N477) );
  INV U1671 ( .IN(N177), .OUT(m1089) );
  NOR2 U1672 ( .A(m1283), .B(m1090), .OUT(N476) );
  INV U1673 ( .IN(N176), .OUT(m1090) );
  NOR2 U1674 ( .A(m1283), .B(m1091), .OUT(N475) );
  INV U1675 ( .IN(N175), .OUT(m1091) );
  NOR2 U1676 ( .A(m1283), .B(m1092), .OUT(N474) );
  INV U1677 ( .IN(N174), .OUT(m1092) );
  NOR2 U1678 ( .A(m1283), .B(m1093), .OUT(N473) );
  INV U1679 ( .IN(N173), .OUT(m1093) );
  NOR2 U1680 ( .A(m1283), .B(m1094), .OUT(N472) );
  INV U1681 ( .IN(N172), .OUT(m1094) );
  NOR2 U1682 ( .A(m1283), .B(m1095), .OUT(N471) );
  INV U1683 ( .IN(N171), .OUT(m1095) );
  NOR2 U1684 ( .A(m1284), .B(m1096), .OUT(N470) );
  INV U1685 ( .IN(N170), .OUT(m1096) );
  NOR2 U1686 ( .A(m1284), .B(m1097), .OUT(N469) );
  INV U1687 ( .IN(N169), .OUT(m1097) );
  NOR2 U1688 ( .A(m1284), .B(m1098), .OUT(N468) );
  INV U1689 ( .IN(N168), .OUT(m1098) );
  NOR2 U1690 ( .A(m1284), .B(m1099), .OUT(N467) );
  INV U1691 ( .IN(N167), .OUT(m1099) );
  NOR2 U1692 ( .A(m1284), .B(m1100), .OUT(N466) );
  INV U1693 ( .IN(N166), .OUT(m1100) );
  NOR2 U1694 ( .A(m1284), .B(m1101), .OUT(N465) );
  INV U1695 ( .IN(N165), .OUT(m1101) );
  NOR2 U1696 ( .A(m1284), .B(m1102), .OUT(N464) );
  INV U1697 ( .IN(N164), .OUT(m1102) );
  NOR2 U1698 ( .A(m1284), .B(m1103), .OUT(N463) );
  INV U1699 ( .IN(N163), .OUT(m1103) );
  NOR2 U1700 ( .A(m1284), .B(m1104), .OUT(N462) );
  INV U1701 ( .IN(N162), .OUT(m1104) );
  NOR2 U1702 ( .A(m1284), .B(m1105), .OUT(N461) );
  INV U1703 ( .IN(N161), .OUT(m1105) );
  NOR2 U1704 ( .A(m1284), .B(m1106), .OUT(N460) );
  INV U1705 ( .IN(N160), .OUT(m1106) );
  NOR2 U1706 ( .A(m1284), .B(m1107), .OUT(N459) );
  INV U1707 ( .IN(N159), .OUT(m1107) );
  NOR2 U1708 ( .A(m1284), .B(m1108), .OUT(N458) );
  INV U1709 ( .IN(N158), .OUT(m1108) );
  NOR2 U1710 ( .A(m1285), .B(m1109), .OUT(N457) );
  INV U1711 ( .IN(N157), .OUT(m1109) );
  NOR2 U1712 ( .A(m1285), .B(m1110), .OUT(N456) );
  INV U1713 ( .IN(N156), .OUT(m1110) );
  NOR2 U1714 ( .A(m1285), .B(m1111), .OUT(N455) );
  INV U1715 ( .IN(N155), .OUT(m1111) );
  NOR2 U1716 ( .A(m1285), .B(m1112), .OUT(N454) );
  INV U1717 ( .IN(N154), .OUT(m1112) );
  NOR2 U1718 ( .A(m1285), .B(m1113), .OUT(N453) );
  INV U1719 ( .IN(N153), .OUT(m1113) );
  NOR2 U1720 ( .A(m1285), .B(m1114), .OUT(N452) );
  INV U1721 ( .IN(N152), .OUT(m1114) );
  NOR2 U1722 ( .A(m1285), .B(m1115), .OUT(N451) );
  INV U1723 ( .IN(N151), .OUT(m1115) );
  NOR2 U1724 ( .A(m1285), .B(m1116), .OUT(N450) );
  INV U1725 ( .IN(N150), .OUT(m1116) );
  NOR2 U1726 ( .A(m1285), .B(m1117), .OUT(N449) );
  INV U1727 ( .IN(N149), .OUT(m1117) );
  NOR2 U1728 ( .A(m1285), .B(m1118), .OUT(N448) );
  INV U1729 ( .IN(N148), .OUT(m1118) );
  NOR2 U1744 ( .A(m1286), .B(m1126), .OUT(N440) );
  INV U1745 ( .IN(N140), .OUT(m1126) );
  NOR2 U1746 ( .A(m1286), .B(m1127), .OUT(N439) );
  INV U1747 ( .IN(N139), .OUT(m1127) );
  NOR2 U1748 ( .A(m1286), .B(m1128), .OUT(N438) );
  INV U1749 ( .IN(N138), .OUT(m1128) );
  NOR2 U1750 ( .A(m1286), .B(m1129), .OUT(N437) );
  INV U1751 ( .IN(N137), .OUT(m1129) );
  NOR2 U1752 ( .A(m1286), .B(m1130), .OUT(N436) );
  INV U1753 ( .IN(N136), .OUT(m1130) );
  NOR2 U1754 ( .A(m1286), .B(m1131), .OUT(N435) );
  INV U1755 ( .IN(N135), .OUT(m1131) );
  NOR2 U1756 ( .A(m1286), .B(m1132), .OUT(N434) );
  INV U1757 ( .IN(N134), .OUT(m1132) );
  NOR2 U1758 ( .A(m1286), .B(m1133), .OUT(N433) );
  INV U1759 ( .IN(N133), .OUT(m1133) );
  NOR2 U1760 ( .A(m1286), .B(m1134), .OUT(N432) );
  INV U1761 ( .IN(N132), .OUT(m1134) );
  NOR2 U1762 ( .A(m1287), .B(m1135), .OUT(N431) );
  INV U1763 ( .IN(N131), .OUT(m1135) );
  NOR2 U1764 ( .A(m1287), .B(m1136), .OUT(N430) );
  INV U1765 ( .IN(N130), .OUT(m1136) );
  NOR2 U1766 ( .A(m1287), .B(m1137), .OUT(N429) );
  INV U1767 ( .IN(N129), .OUT(m1137) );
  NOR2 U1768 ( .A(m1287), .B(m1138), .OUT(N428) );
  INV U1769 ( .IN(N128), .OUT(m1138) );
  NOR2 U1786 ( .A(m1287), .B(m1147), .OUT(N419) );
  INV U1787 ( .IN(N119), .OUT(m1147) );
  NOR2 U1788 ( .A(m1287), .B(m1148), .OUT(N418) );
  INV U1789 ( .IN(N118), .OUT(m1148) );
  NOR2 U1790 ( .A(m1287), .B(m1149), .OUT(N417) );
  INV U1791 ( .IN(N117), .OUT(m1149) );
  NOR2 U1792 ( .A(m1287), .B(m1150), .OUT(N416) );
  INV U1793 ( .IN(N116), .OUT(m1150) );
  NOR2 U1794 ( .A(m1287), .B(m1151), .OUT(N415) );
  INV U1795 ( .IN(N115), .OUT(m1151) );
  NOR2 U1796 ( .A(m1287), .B(m1152), .OUT(N414) );
  INV U1797 ( .IN(N114), .OUT(m1152) );
  NOR2 U1798 ( .A(m1287), .B(m1153), .OUT(N413) );
  INV U1799 ( .IN(N113), .OUT(m1153) );
  NOR2 U1800 ( .A(m1287), .B(m1154), .OUT(N412) );
  INV U1801 ( .IN(N112), .OUT(m1154) );
  NOR2 U1802 ( .A(m1287), .B(m1155), .OUT(N411) );
  INV U1803 ( .IN(N111), .OUT(m1155) );
  NOR2 U1804 ( .A(m1288), .B(m1156), .OUT(N410) );
  INV U1805 ( .IN(N110), .OUT(m1156) );
  NOR2 U1806 ( .A(m1288), .B(m1157), .OUT(N409) );
  INV U1807 ( .IN(N109), .OUT(m1157) );
  NOR2 U1808 ( .A(m1288), .B(m1158), .OUT(N408) );
  INV U1809 ( .IN(N108), .OUT(m1158) );
  NOR2 U1810 ( .A(m1288), .B(m1159), .OUT(N407) );
  INV U1811 ( .IN(acc[19]), .OUT(m1159) );
  NOR2 U1812 ( .A(m1288), .B(m1160), .OUT(N406) );
  INV U1813 ( .IN(acc[18]), .OUT(m1160) );
  NOR2 U1814 ( .A(m1288), .B(m1161), .OUT(N405) );
  INV U1815 ( .IN(acc[17]), .OUT(m1161) );
  NOR2 U1816 ( .A(m1288), .B(m1162), .OUT(N404) );
  INV U1817 ( .IN(acc[16]), .OUT(m1162) );
  NOR2 U1818 ( .A(m1288), .B(m1163), .OUT(N403) );
  INV U1819 ( .IN(acc[15]), .OUT(m1163) );
  NOR2 U1820 ( .A(m1288), .B(m1164), .OUT(N402) );
  INV U1821 ( .IN(acc[14]), .OUT(m1164) );
  NOR2 U1822 ( .A(m1288), .B(m1165), .OUT(N401) );
  INV U1823 ( .IN(acc[13]), .OUT(m1165) );
  NOR2 U1824 ( .A(m1288), .B(m1166), .OUT(N400) );
  INV U1825 ( .IN(acc[12]), .OUT(m1166) );
  NOR2 U1826 ( .A(m1288), .B(m1167), .OUT(N399) );
  INV U1827 ( .IN(acc[11]), .OUT(m1167) );
  NOR2 U1828 ( .A(m1288), .B(m1168), .OUT(N398) );
  INV U1829 ( .IN(acc[10]), .OUT(m1168) );
  NOR2 U1830 ( .A(m1289), .B(m1169), .OUT(N397) );
  INV U1831 ( .IN(acc[9]), .OUT(m1169) );
  NOR2 U1832 ( .A(m1289), .B(m1170), .OUT(N396) );
  INV U1833 ( .IN(acc[8]), .OUT(m1170) );
  NOR2 U1834 ( .A(m1289), .B(m1171), .OUT(N395) );
  INV U1835 ( .IN(acc[7]), .OUT(m1171) );
  NOR2 U1836 ( .A(m1289), .B(m1172), .OUT(N394) );
  INV U1837 ( .IN(acc[6]), .OUT(m1172) );
  NOR2 U1838 ( .A(m1289), .B(m1173), .OUT(N393) );
  INV U1839 ( .IN(acc[5]), .OUT(m1173) );
  NOR2 U1840 ( .A(m1289), .B(m1174), .OUT(N392) );
  INV U1841 ( .IN(acc[4]), .OUT(m1174) );
  NOR2 U1842 ( .A(m1289), .B(m1175), .OUT(N391) );
  INV U1843 ( .IN(acc[3]), .OUT(m1175) );
  NOR2 U1844 ( .A(m1289), .B(m1176), .OUT(N390) );
  INV U1845 ( .IN(acc[2]), .OUT(m1176) );
  NOR2 U1846 ( .A(m1289), .B(m1177), .OUT(N389) );
  INV U1847 ( .IN(acc[1]), .OUT(m1177) );
  NOR2 U1848 ( .A(m1289), .B(m1178), .OUT(N388) );
  INV U1849 ( .IN(acc[0]), .OUT(m1178) );
  INV \mult_83/AN1_7  ( .IN(\Samples[12][7] ), .OUT(\mult_83/A_not[7] ) );
  INV \mult_83/AN1_6  ( .IN(\Samples[12][6] ), .OUT(\mult_83/A_notx [6]) );
  INV \mult_83/AN1_5  ( .IN(\Samples[12][5] ), .OUT(\mult_83/A_notx [5]) );
  INV \mult_83/AN1_4  ( .IN(\Samples[12][4] ), .OUT(\mult_83/A_notx [4]) );
  INV \mult_83/AN1_3  ( .IN(\Samples[12][3] ), .OUT(\mult_83/A_notx [3]) );
  INV \mult_83/AN1_2  ( .IN(\Samples[12][2] ), .OUT(\mult_83/A_notx [2]) );
  INV \mult_83/AN1_1  ( .IN(\Samples[12][1] ), .OUT(\mult_83/A_notx [1]) );
  INV \mult_83/AN1_0  ( .IN(\Samples[12][0] ), .OUT(\mult_83/A_notx [0]) );
  XOR2 \mult_80/FS_1/U3_C_0_2_0  ( .A(\mult_80/FS_1/PG_int[0][2][0] ), .B(
        \mult_80/FS_1/C[1][2][0] ), .OUT(N83) );
  NAND2 \mult_80/FS_1/U3_B_0_1_3  ( .A(\mult_80/FS_1/G_n_int[0][1][3] ), .B(
        \mult_80/FS_1/P[0][1][3] ), .OUT(m2576) );
  NAND2 \mult_80/FS_1/U2_0_1_3  ( .A(\mult_80/A1[7] ), .B(\mult_80/A2[7] ), 
        .OUT(\mult_80/FS_1/G_n_int[0][1][3] ) );
  NAND2 \mult_80/FS_1/U1_0_1_3  ( .A(m2574), .B(m2575), .OUT(
        \mult_80/FS_1/P[0][1][3] ) );
  INV \mult_80/AN1_7  ( .IN(\Samples[9][7] ), .OUT(\mult_80/A_not[7] ) );
  INV \mult_80/AN1_6  ( .IN(\Samples[9][6] ), .OUT(\mult_80/A_notx [6]) );
  INV \mult_80/AN1_5  ( .IN(\Samples[9][5] ), .OUT(\mult_80/A_notx [5]) );
  INV \mult_80/AN1_4  ( .IN(\Samples[9][4] ), .OUT(\mult_80/A_notx [4]) );
  INV \mult_80/AN1_3  ( .IN(\Samples[9][3] ), .OUT(\mult_80/A_notx [3]) );
  INV \mult_80/AN1_2  ( .IN(\Samples[9][2] ), .OUT(\mult_80/A_notx [2]) );
  INV \mult_80/AN1_1  ( .IN(\Samples[9][1] ), .OUT(\mult_80/A_notx [1]) );
  INV \mult_80/AN1_0  ( .IN(\Samples[9][0] ), .OUT(\mult_80/A_notx [0]) );
  INV \mult_77/AN1_7  ( .IN(\Samples[7][7] ), .OUT(\mult_77/A_not[7] ) );
  INV \mult_77/AN1_6  ( .IN(\Samples[7][6] ), .OUT(\mult_77/A_notx [6]) );
  INV \mult_77/AN1_5  ( .IN(\Samples[7][5] ), .OUT(\mult_77/A_notx [5]) );
  INV \mult_77/AN1_4  ( .IN(\Samples[7][4] ), .OUT(\mult_77/A_notx [4]) );
  INV \mult_77/AN1_3  ( .IN(\Samples[7][3] ), .OUT(\mult_77/A_notx [3]) );
  INV \mult_77/AN1_2  ( .IN(\Samples[7][2] ), .OUT(\mult_77/A_notx [2]) );
  INV \mult_77/AN1_1  ( .IN(\Samples[7][1] ), .OUT(\mult_77/A_notx [1]) );
  INV \mult_77/AN1_0  ( .IN(\Samples[7][0] ), .OUT(\mult_77/A_notx [0]) );
  XOR2 \mult_76/FS_1/U3_C_0_2_0  ( .A(\mult_76/FS_1/PG_int[0][2][0] ), .B(
        \mult_76/FS_1/C[1][2][0] ), .OUT(N59) );
  NAND2 \mult_76/FS_1/U3_B_0_1_3  ( .A(\mult_76/FS_1/G_n_int[0][1][3] ), .B(
        \mult_76/FS_1/P[0][1][3] ), .OUT(m2534) );
  NAND2 \mult_76/FS_1/U2_0_1_3  ( .A(\mult_76/A1[7] ), .B(\mult_76/A2[7] ), 
        .OUT(\mult_76/FS_1/G_n_int[0][1][3] ) );
  NAND2 \mult_76/FS_1/U1_0_1_3  ( .A(m2532), .B(m2533), .OUT(
        \mult_76/FS_1/P[0][1][3] ) );
  INV \mult_76/AN1_7  ( .IN(\Samples[6][7] ), .OUT(\mult_76/A_not[7] ) );
  INV \mult_76/AN1_6  ( .IN(\Samples[6][6] ), .OUT(\mult_76/A_notx [6]) );
  INV \mult_76/AN1_5  ( .IN(\Samples[6][5] ), .OUT(\mult_76/A_notx [5]) );
  INV \mult_76/AN1_4  ( .IN(\Samples[6][4] ), .OUT(\mult_76/A_notx [4]) );
  INV \mult_76/AN1_3  ( .IN(\Samples[6][3] ), .OUT(\mult_76/A_notx [3]) );
  INV \mult_76/AN1_2  ( .IN(\Samples[6][2] ), .OUT(\mult_76/A_notx [2]) );
  INV \mult_76/AN1_1  ( .IN(\Samples[6][1] ), .OUT(\mult_76/A_notx [1]) );
  INV \mult_76/AN1_0  ( .IN(\Samples[6][0] ), .OUT(\mult_76/A_notx [0]) );
  XOR2 \mult_74/FS_1/U3_C_0_2_0  ( .A(\mult_74/FS_1/PG_int[0][2][0] ), .B(
        \mult_74/FS_1/C[1][2][0] ), .OUT(N48) );
  NAND2 \mult_74/FS_1/U3_B_0_1_3  ( .A(\mult_74/FS_1/G_n_int[0][1][3] ), .B(
        \mult_74/FS_1/P[0][1][3] ), .OUT(m2513) );
  NAND2 \mult_74/FS_1/U2_0_1_3  ( .A(\mult_74/A1[7] ), .B(\mult_74/A2[7] ), 
        .OUT(\mult_74/FS_1/G_n_int[0][1][3] ) );
  NAND2 \mult_74/FS_1/U1_0_1_3  ( .A(m2511), .B(m2512), .OUT(
        \mult_74/FS_1/P[0][1][3] ) );
  INV \mult_74/AN1_7  ( .IN(\Samples[4][7] ), .OUT(\mult_74/A_not[7] ) );
  INV \mult_74/AN1_6  ( .IN(\Samples[4][6] ), .OUT(\mult_74/A_notx [6]) );
  INV \mult_74/AN1_5  ( .IN(\Samples[4][5] ), .OUT(\mult_74/A_notx [5]) );
  INV \mult_74/AN1_4  ( .IN(\Samples[4][4] ), .OUT(\mult_74/A_notx [4]) );
  INV \mult_74/AN1_3  ( .IN(\Samples[4][3] ), .OUT(\mult_74/A_notx [3]) );
  INV \mult_74/AN1_2  ( .IN(\Samples[4][2] ), .OUT(\mult_74/A_notx [2]) );
  INV \mult_74/AN1_1  ( .IN(\Samples[4][1] ), .OUT(\mult_74/A_notx [1]) );
  INV \mult_74/AN1_0  ( .IN(\Samples[4][0] ), .OUT(\mult_74/A_notx [0]) );
  INV \mult_72/AN1_7  ( .IN(\Samples[2][7] ), .OUT(\mult_72/A_not[7] ) );
  INV \mult_72/AN1_6  ( .IN(\Samples[2][6] ), .OUT(\mult_72/A_notx [6]) );
  INV \mult_72/AN1_5  ( .IN(\Samples[2][5] ), .OUT(\mult_72/A_notx [5]) );
  INV \mult_72/AN1_4  ( .IN(\Samples[2][4] ), .OUT(\mult_72/A_notx [4]) );
  INV \mult_72/AN1_3  ( .IN(\Samples[2][3] ), .OUT(\mult_72/A_notx [3]) );
  INV \mult_72/AN1_2  ( .IN(\Samples[2][2] ), .OUT(\mult_72/A_notx [2]) );
  INV \mult_72/AN1_1  ( .IN(\Samples[2][1] ), .OUT(\mult_72/A_notx [1]) );
  INV \mult_72/AN1_0  ( .IN(\Samples[2][0] ), .OUT(\mult_72/A_notx [0]) );
  XOR2 \mult_71/FS_1/U3_C_0_2_0  ( .A(\mult_71/FS_1/PG_int[0][2][0] ), .B(
        \mult_71/FS_1/C[1][2][0] ), .OUT(N24) );
  NAND2 \mult_71/FS_1/U3_B_0_1_3  ( .A(\mult_71/FS_1/G_n_int[0][1][3] ), .B(
        \mult_71/FS_1/P[0][1][3] ), .OUT(m2471) );
  NAND2 \mult_71/FS_1/U2_0_1_3  ( .A(\mult_71/A1[7] ), .B(\mult_71/A2[7] ), 
        .OUT(\mult_71/FS_1/G_n_int[0][1][3] ) );
  NAND2 \mult_71/FS_1/U1_0_1_3  ( .A(m2469), .B(m2470), .OUT(
        \mult_71/FS_1/P[0][1][3] ) );
  INV \mult_71/AN1_7  ( .IN(\Samples[1][7] ), .OUT(\mult_71/A_not[7] ) );
  INV \mult_71/AN1_6  ( .IN(\Samples[1][6] ), .OUT(\mult_71/A_notx [6]) );
  INV \mult_71/AN1_5  ( .IN(\Samples[1][5] ), .OUT(\mult_71/A_notx [5]) );
  INV \mult_71/AN1_4  ( .IN(\Samples[1][4] ), .OUT(\mult_71/A_notx [4]) );
  INV \mult_71/AN1_3  ( .IN(\Samples[1][3] ), .OUT(\mult_71/A_notx [3]) );
  INV \mult_71/AN1_2  ( .IN(\Samples[1][2] ), .OUT(\mult_71/A_notx [2]) );
  INV \mult_71/AN1_1  ( .IN(\Samples[1][1] ), .OUT(\mult_71/A_notx [1]) );
  INV \mult_71/AN1_0  ( .IN(\Samples[1][0] ), .OUT(\mult_71/A_notx [0]) );
  XOR2 \mult_69/FS_1/U3_C_0_2_0  ( .A(\mult_69/FS_1/PG_int[0][2][0] ), .B(
        \mult_69/FS_1/C[1][2][0] ), .OUT(N13) );
  NAND2 \mult_69/FS_1/U3_B_0_1_3  ( .A(\mult_69/FS_1/G_n_int[0][1][3] ), .B(
        \mult_69/FS_1/P[0][1][3] ), .OUT(m2450) );
  NAND2 \mult_69/FS_1/U2_0_1_3  ( .A(\mult_69/A1[7] ), .B(\mult_69/A2[7] ), 
        .OUT(\mult_69/FS_1/G_n_int[0][1][3] ) );
  NAND2 \mult_69/FS_1/U1_0_1_3  ( .A(m2448), .B(m2449), .OUT(
        \mult_69/FS_1/P[0][1][3] ) );
  INV \mult_69/AN1_7  ( .IN(Data_in[7]), .OUT(\mult_69/A_not[7] ) );
  INV \mult_69/AN1_6  ( .IN(Data_in[6]), .OUT(\mult_69/A_notx [6]) );
  INV \mult_69/AN1_5  ( .IN(Data_in[5]), .OUT(\mult_69/A_notx [5]) );
  INV \mult_69/AN1_4  ( .IN(Data_in[4]), .OUT(\mult_69/A_notx [4]) );
  INV \mult_69/AN1_3  ( .IN(Data_in[3]), .OUT(\mult_69/A_notx [3]) );
  INV \mult_69/AN1_2  ( .IN(Data_in[2]), .OUT(\mult_69/A_notx [2]) );
  INV \mult_69/AN1_1  ( .IN(Data_in[1]), .OUT(\mult_69/A_notx [1]) );
  INV \mult_69/AN1_0  ( .IN(Data_in[0]), .OUT(\mult_69/A_notx [0]) );
  XOR2 \mult_82/FS_1/U3_C_0_2_0  ( .A(\mult_82/FS_1/PG_int[0][2][0] ), .B(
        \mult_82/FS_1/C[1][2][0] ), .OUT(N94) );
  NAND2 \mult_82/FS_1/U3_B_0_1_3  ( .A(\mult_82/FS_1/G_n_int[0][1][3] ), .B(
        \mult_82/FS_1/P[0][1][3] ), .OUT(m2428) );
  NAND2 \mult_82/FS_1/U2_0_1_3  ( .A(\mult_82/A1[7] ), .B(\mult_82/A2[7] ), 
        .OUT(\mult_82/FS_1/G_n_int[0][1][3] ) );
  NAND2 \mult_82/FS_1/U1_0_1_3  ( .A(m2426), .B(m2427), .OUT(
        \mult_82/FS_1/P[0][1][3] ) );
  INV \mult_82/AN1_7  ( .IN(\Samples[11][7] ), .OUT(\mult_82/A_not[7] ) );
  INV \mult_82/AN1_6  ( .IN(\Samples[11][6] ), .OUT(\mult_82/A_notx [6]) );
  INV \mult_82/AN1_5  ( .IN(\Samples[11][5] ), .OUT(\mult_82/A_notx [5]) );
  INV \mult_82/AN1_4  ( .IN(\Samples[11][4] ), .OUT(\mult_82/A_notx [4]) );
  INV \mult_82/AN1_3  ( .IN(\Samples[11][3] ), .OUT(\mult_82/A_notx [3]) );
  INV \mult_82/AN1_2  ( .IN(\Samples[11][2] ), .OUT(\mult_82/A_notx [2]) );
  INV \mult_82/AN1_1  ( .IN(\Samples[11][1] ), .OUT(\mult_82/A_notx [1]) );
  INV \mult_82/AN1_0  ( .IN(\Samples[11][0] ), .OUT(\mult_82/A_notx [0]) );
  XOR2 U1850 ( .A(1'b1), .B(m2118), .OUT(N349) );
  XOR2 U1851 ( .A(1'b1), .B(\PR_add[11][1] ), .OUT(m2118) );
  XOR2 U1852 ( .A(1'b1), .B(m2143), .OUT(N249) );
  XOR2 U1853 ( .A(1'b1), .B(\PR_add[6][1] ), .OUT(m2143) );
  XOR2 U1854 ( .A(1'b1), .B(m2168), .OUT(N149) );
  XOR2 U1855 ( .A(1'b1), .B(\PR_add[1][1] ), .OUT(m2168) );
  NAND2 U1856 ( .A(\PR_mul[3][2] ), .B(\PR_add[1][2] ), .OUT(m1923) );
  NAND2 U1857 ( .A(\PR_mul[8][2] ), .B(\PR_add[6][2] ), .OUT(m1843) );
  NAND2 U1858 ( .A(\PR_mul[13][2] ), .B(\PR_add[11][2] ), .OUT(m1763) );
  INV U1860 ( .IN(m1187), .OUT(m1180) );
  INV U1861 ( .IN(m1187), .OUT(m1181) );
  INV U1862 ( .IN(m1187), .OUT(m1182) );
  INV U1863 ( .IN(m1186), .OUT(m1183) );
  INV U1864 ( .IN(m1186), .OUT(m1184) );
  INV U1865 ( .IN(m1186), .OUT(m1185) );
  INV U1866 ( .IN(m631), .OUT(m1186) );
  INV U1867 ( .IN(m631), .OUT(m1187) );
  INV U1868 ( .IN(m1251), .OUT(m1188) );
  INV U1869 ( .IN(m1251), .OUT(m1189) );
  INV U1870 ( .IN(m1251), .OUT(m1190) );
  INV U1871 ( .IN(m1250), .OUT(m1191) );
  INV U1872 ( .IN(m1250), .OUT(m1192) );
  INV U1873 ( .IN(m1250), .OUT(m1193) );
  INV U1874 ( .IN(m1249), .OUT(m1194) );
  INV U1875 ( .IN(m1249), .OUT(m1195) );
  INV U1876 ( .IN(m1249), .OUT(m1196) );
  INV U1877 ( .IN(m1248), .OUT(m1197) );
  INV U1878 ( .IN(m1248), .OUT(m1198) );
  INV U1879 ( .IN(m1248), .OUT(m1199) );
  INV U1880 ( .IN(m1247), .OUT(m1200) );
  INV U1881 ( .IN(m1247), .OUT(m1201) );
  INV U1882 ( .IN(m1247), .OUT(m1202) );
  INV U1883 ( .IN(m1246), .OUT(m1203) );
  INV U1884 ( .IN(m1246), .OUT(m1204) );
  INV U1885 ( .IN(m1246), .OUT(m1205) );
  INV U1886 ( .IN(m1245), .OUT(m1206) );
  INV U1887 ( .IN(m1245), .OUT(m1207) );
  INV U1888 ( .IN(m1245), .OUT(m1208) );
  INV U1889 ( .IN(m1244), .OUT(m1209) );
  INV U1890 ( .IN(m1244), .OUT(m1210) );
  INV U1891 ( .IN(m1244), .OUT(m1211) );
  INV U1892 ( .IN(m1243), .OUT(m1212) );
  INV U1893 ( .IN(m1243), .OUT(m1213) );
  INV U1894 ( .IN(m1243), .OUT(m1214) );
  INV U1895 ( .IN(m1242), .OUT(m1215) );
  INV U1896 ( .IN(m1242), .OUT(m1216) );
  INV U1897 ( .IN(m1242), .OUT(m1217) );
  INV U1898 ( .IN(m1241), .OUT(m1218) );
  INV U1899 ( .IN(m1241), .OUT(m1219) );
  INV U1900 ( .IN(m1241), .OUT(m1220) );
  INV U1901 ( .IN(m1240), .OUT(m1221) );
  INV U1902 ( .IN(m1240), .OUT(m1222) );
  INV U1903 ( .IN(m1240), .OUT(m1223) );
  INV U1904 ( .IN(m1239), .OUT(m1224) );
  INV U1905 ( .IN(m1239), .OUT(m1225) );
  INV U1906 ( .IN(m1239), .OUT(m1226) );
  INV U1907 ( .IN(m1238), .OUT(m1227) );
  INV U1908 ( .IN(m1238), .OUT(m1228) );
  INV U1909 ( .IN(m1238), .OUT(m1229) );
  INV U1910 ( .IN(m1237), .OUT(m1230) );
  INV U1911 ( .IN(m1237), .OUT(m1231) );
  INV U1912 ( .IN(m1237), .OUT(m1232) );
  INV U1913 ( .IN(m1236), .OUT(m1233) );
  INV U1914 ( .IN(m1236), .OUT(m1234) );
  INV U1915 ( .IN(m1236), .OUT(m1235) );
  INV U1916 ( .IN(m1180), .OUT(m1236) );
  INV U1917 ( .IN(m1180), .OUT(m1237) );
  INV U1918 ( .IN(m1180), .OUT(m1238) );
  INV U1919 ( .IN(m1181), .OUT(m1239) );
  INV U1920 ( .IN(m1181), .OUT(m1240) );
  INV U1921 ( .IN(m1181), .OUT(m1241) );
  INV U1922 ( .IN(m1182), .OUT(m1242) );
  INV U1923 ( .IN(m1182), .OUT(m1243) );
  INV U1924 ( .IN(m1182), .OUT(m1244) );
  INV U1925 ( .IN(m1183), .OUT(m1245) );
  INV U1926 ( .IN(m1183), .OUT(m1246) );
  INV U1927 ( .IN(m1183), .OUT(m1247) );
  INV U1928 ( .IN(m1184), .OUT(m1248) );
  INV U1929 ( .IN(m1184), .OUT(m1249) );
  INV U1930 ( .IN(m1184), .OUT(m1250) );
  INV U1931 ( .IN(m1185), .OUT(m1251) );
  INV U1932 ( .IN(m1302), .OUT(m1252) );
  INV U1933 ( .IN(m1302), .OUT(m1253) );
  INV U1934 ( .IN(m1301), .OUT(m1254) );
  INV U1935 ( .IN(m1301), .OUT(m1255) );
  INV U1936 ( .IN(m1301), .OUT(m1256) );
  INV U1937 ( .IN(m1300), .OUT(m1257) );
  INV U1938 ( .IN(m1300), .OUT(m1258) );
  INV U1939 ( .IN(m1300), .OUT(m1259) );
  INV U1940 ( .IN(m1299), .OUT(m1260) );
  INV U1941 ( .IN(m1299), .OUT(m1261) );
  INV U1942 ( .IN(m1299), .OUT(m1262) );
  INV U1943 ( .IN(m1298), .OUT(m1263) );
  INV U1944 ( .IN(m1298), .OUT(m1264) );
  INV U1945 ( .IN(m1298), .OUT(m1265) );
  INV U1946 ( .IN(m1297), .OUT(m1266) );
  INV U1947 ( .IN(m1297), .OUT(m1267) );
  INV U1948 ( .IN(m1297), .OUT(m1268) );
  INV U1949 ( .IN(m1296), .OUT(m1269) );
  INV U1950 ( .IN(m1296), .OUT(m1270) );
  INV U1951 ( .IN(m1296), .OUT(m1271) );
  INV U1952 ( .IN(m1295), .OUT(m1272) );
  INV U1953 ( .IN(m1295), .OUT(m1273) );
  INV U1954 ( .IN(m1295), .OUT(m1274) );
  INV U1955 ( .IN(m1294), .OUT(m1275) );
  INV U1956 ( .IN(m1294), .OUT(m1276) );
  INV U1957 ( .IN(m1294), .OUT(m1277) );
  INV U1958 ( .IN(m1293), .OUT(m1278) );
  INV U1959 ( .IN(m1293), .OUT(m1279) );
  INV U1960 ( .IN(m1293), .OUT(m1280) );
  INV U1961 ( .IN(m1292), .OUT(m1281) );
  INV U1962 ( .IN(m1292), .OUT(m1282) );
  INV U1963 ( .IN(m1292), .OUT(m1283) );
  INV U1964 ( .IN(m1291), .OUT(m1284) );
  INV U1965 ( .IN(m1291), .OUT(m1285) );
  INV U1966 ( .IN(m1291), .OUT(m1286) );
  INV U1967 ( .IN(m1290), .OUT(m1287) );
  INV U1968 ( .IN(m1290), .OUT(m1288) );
  INV U1969 ( .IN(m1290), .OUT(m1289) );
  INV U1970 ( .IN(reset), .OUT(m1290) );
  INV U1971 ( .IN(reset), .OUT(m1291) );
  INV U1972 ( .IN(reset), .OUT(m1292) );
  INV U1973 ( .IN(reset), .OUT(m1293) );
  INV U1974 ( .IN(reset), .OUT(m1294) );
  INV U1975 ( .IN(reset), .OUT(m1295) );
  INV U1976 ( .IN(reset), .OUT(m1296) );
  INV U1977 ( .IN(reset), .OUT(m1297) );
  INV U1978 ( .IN(reset), .OUT(m1298) );
  INV U1979 ( .IN(reset), .OUT(m1299) );
  INV U1980 ( .IN(reset), .OUT(m1300) );
  INV U1981 ( .IN(reset), .OUT(m1301) );
  INV U1982 ( .IN(reset), .OUT(m1302) );
  INV U1983 ( .IN(reset), .OUT(m1303) );
  INV U1984 ( .IN(reset), .OUT(m1304) );
  INV U1985 ( .IN(reset), .OUT(m1305) );
  INV U1986 ( .IN(reset), .OUT(m1306) );
  INV U1987 ( .IN(reset), .OUT(m1307) );
  INV U1988 ( .IN(reset), .OUT(m1308) );
  INV U1989 ( .IN(reset), .OUT(m1309) );
  INV U1990 ( .IN(reset), .OUT(m1310) );
  INV U1991 ( .IN(reset), .OUT(m1311) );
  INV U1992 ( .IN(reset), .OUT(m1312) );
  INV U1993 ( .IN(reset), .OUT(m1313) );
  INV U1994 ( .IN(reset), .OUT(m1314) );
  INV U1995 ( .IN(reset), .OUT(m1315) );
  INV U2002 ( .IN(m2412), .OUT(\mult_82/FS_1/TEMP_P[0][0][0] ) );
  INV U2003 ( .IN(m2434), .OUT(\mult_69/FS_1/TEMP_P[0][0][0] ) );
  INV U2004 ( .IN(m2455), .OUT(\mult_71/FS_1/TEMP_P[0][0][0] ) );
  INV U2005 ( .IN(m2477), .OUT(\mult_72/FS_1/TEMP_P[0][0][0] ) );
  INV U2006 ( .IN(m2497), .OUT(\mult_74/FS_1/TEMP_P[0][0][0] ) );
  INV U2007 ( .IN(m2518), .OUT(\mult_76/FS_1/TEMP_P[0][0][0] ) );
  INV U2008 ( .IN(m2540), .OUT(\mult_77/FS_1/TEMP_P[0][0][0] ) );
  INV U2009 ( .IN(m2560), .OUT(\mult_80/FS_1/TEMP_P[0][0][0] ) );
  INV U2010 ( .IN(m2581), .OUT(\mult_83/FS_1/TEMP_P[0][0][0] ) );
  INV U2011 ( .IN(\mult_83/FS_1/TEMP_P[0][0][0] ), .OUT(m2582) );
  INV U2012 ( .IN(m2583), .OUT(\mult_83/FS_1/P[0][0][1] ) );
  INV U2013 ( .IN(\mult_82/FS_1/TEMP_P[0][0][0] ), .OUT(m2413) );
  INV U2014 ( .IN(m2414), .OUT(\mult_82/FS_1/P[0][0][1] ) );
  INV U2015 ( .IN(\mult_80/FS_1/TEMP_P[0][0][0] ), .OUT(m2561) );
  INV U2016 ( .IN(m2562), .OUT(\mult_80/FS_1/P[0][0][1] ) );
  INV U2017 ( .IN(\mult_77/FS_1/TEMP_P[0][0][0] ), .OUT(m2541) );
  INV U2018 ( .IN(m2542), .OUT(\mult_77/FS_1/P[0][0][1] ) );
  INV U2019 ( .IN(\mult_76/FS_1/TEMP_P[0][0][0] ), .OUT(m2519) );
  INV U2020 ( .IN(m2520), .OUT(\mult_76/FS_1/P[0][0][1] ) );
  INV U2021 ( .IN(\mult_74/FS_1/TEMP_P[0][0][0] ), .OUT(m2498) );
  INV U2022 ( .IN(m2499), .OUT(\mult_74/FS_1/P[0][0][1] ) );
  INV U2023 ( .IN(\mult_72/FS_1/TEMP_P[0][0][0] ), .OUT(m2478) );
  INV U2024 ( .IN(m2479), .OUT(\mult_72/FS_1/P[0][0][1] ) );
  INV U2025 ( .IN(\mult_71/FS_1/TEMP_P[0][0][0] ), .OUT(m2456) );
  INV U2026 ( .IN(m2457), .OUT(\mult_71/FS_1/P[0][0][1] ) );
  INV U2027 ( .IN(\mult_83/FS_1/P[0][0][1] ), .OUT(m2584) );
  INV U2028 ( .IN(m2585), .OUT(\mult_83/FS_1/P[0][0][2] ) );
  INV U2029 ( .IN(\mult_82/FS_1/P[0][0][1] ), .OUT(m2415) );
  INV U2030 ( .IN(m2416), .OUT(\mult_82/FS_1/P[0][0][2] ) );
  INV U2031 ( .IN(\mult_80/FS_1/P[0][0][1] ), .OUT(m2563) );
  INV U2032 ( .IN(m2564), .OUT(\mult_80/FS_1/P[0][0][2] ) );
  INV U2033 ( .IN(\mult_77/FS_1/P[0][0][1] ), .OUT(m2543) );
  INV U2034 ( .IN(m2544), .OUT(\mult_77/FS_1/P[0][0][2] ) );
  INV U2035 ( .IN(\mult_76/FS_1/P[0][0][1] ), .OUT(m2521) );
  INV U2036 ( .IN(m2522), .OUT(\mult_76/FS_1/P[0][0][2] ) );
  INV U2037 ( .IN(\mult_74/FS_1/P[0][0][1] ), .OUT(m2500) );
  INV U2038 ( .IN(m2501), .OUT(\mult_74/FS_1/P[0][0][2] ) );
  INV U2039 ( .IN(\mult_72/FS_1/P[0][0][1] ), .OUT(m2480) );
  INV U2040 ( .IN(m2481), .OUT(\mult_72/FS_1/P[0][0][2] ) );
  INV U2041 ( .IN(\mult_71/FS_1/P[0][0][1] ), .OUT(m2458) );
  INV U2042 ( .IN(m2459), .OUT(\mult_71/FS_1/P[0][0][2] ) );
  INV U2043 ( .IN(\mult_83/FS_1/P[0][0][2] ), .OUT(m2586) );
  INV U2044 ( .IN(m2587), .OUT(\mult_83/FS_1/P[0][0][3] ) );
  INV U2045 ( .IN(\mult_82/FS_1/P[0][0][2] ), .OUT(m2417) );
  INV U2046 ( .IN(m2418), .OUT(\mult_82/FS_1/P[0][0][3] ) );
  INV U2047 ( .IN(\mult_80/FS_1/P[0][0][2] ), .OUT(m2565) );
  INV U2048 ( .IN(m2566), .OUT(\mult_80/FS_1/P[0][0][3] ) );
  INV U2049 ( .IN(\mult_77/FS_1/P[0][0][2] ), .OUT(m2545) );
  INV U2050 ( .IN(m2546), .OUT(\mult_77/FS_1/P[0][0][3] ) );
  INV U2051 ( .IN(\mult_76/FS_1/P[0][0][2] ), .OUT(m2523) );
  INV U2052 ( .IN(m2524), .OUT(\mult_76/FS_1/P[0][0][3] ) );
  INV U2053 ( .IN(\mult_74/FS_1/P[0][0][2] ), .OUT(m2502) );
  INV U2054 ( .IN(m2503), .OUT(\mult_74/FS_1/P[0][0][3] ) );
  INV U2055 ( .IN(\mult_72/FS_1/P[0][0][2] ), .OUT(m2482) );
  INV U2056 ( .IN(m2483), .OUT(\mult_72/FS_1/P[0][0][3] ) );
  INV U2057 ( .IN(\mult_71/FS_1/P[0][0][2] ), .OUT(m2460) );
  INV U2058 ( .IN(m2461), .OUT(\mult_71/FS_1/P[0][0][3] ) );
  INV U2059 ( .IN(\mult_83/FS_1/P[0][0][3] ), .OUT(m2588) );
  INV U2060 ( .IN(m2589), .OUT(\mult_83/FS_1/TEMP_P[0][1][0] ) );
  INV U2061 ( .IN(\mult_82/FS_1/P[0][0][3] ), .OUT(m2419) );
  INV U2062 ( .IN(m2420), .OUT(\mult_82/FS_1/TEMP_P[0][1][0] ) );
  INV U2063 ( .IN(\mult_80/FS_1/P[0][0][3] ), .OUT(m2567) );
  INV U2064 ( .IN(m2568), .OUT(\mult_80/FS_1/TEMP_P[0][1][0] ) );
  INV U2065 ( .IN(\mult_77/FS_1/P[0][0][3] ), .OUT(m2547) );
  INV U2066 ( .IN(m2548), .OUT(\mult_77/FS_1/TEMP_P[0][1][0] ) );
  INV U2067 ( .IN(\mult_76/FS_1/P[0][0][3] ), .OUT(m2525) );
  INV U2068 ( .IN(m2526), .OUT(\mult_76/FS_1/TEMP_P[0][1][0] ) );
  INV U2069 ( .IN(\mult_74/FS_1/P[0][0][3] ), .OUT(m2504) );
  INV U2070 ( .IN(m2505), .OUT(\mult_74/FS_1/TEMP_P[0][1][0] ) );
  INV U2071 ( .IN(\mult_72/FS_1/P[0][0][3] ), .OUT(m2484) );
  INV U2072 ( .IN(m2485), .OUT(\mult_72/FS_1/TEMP_P[0][1][0] ) );
  INV U2073 ( .IN(\mult_71/FS_1/P[0][0][3] ), .OUT(m2462) );
  INV U2074 ( .IN(m2463), .OUT(\mult_71/FS_1/TEMP_P[0][1][0] ) );
  INV U2075 ( .IN(\mult_83/FS_1/TEMP_P[0][1][0] ), .OUT(m2590) );
  INV U2076 ( .IN(m2591), .OUT(\mult_83/FS_1/P[0][1][1] ) );
  INV U2077 ( .IN(\mult_82/FS_1/TEMP_P[0][1][0] ), .OUT(m2421) );
  INV U2078 ( .IN(m2422), .OUT(\mult_82/FS_1/P[0][1][1] ) );
  INV U2079 ( .IN(\mult_80/FS_1/TEMP_P[0][1][0] ), .OUT(m2569) );
  INV U2080 ( .IN(m2570), .OUT(\mult_80/FS_1/P[0][1][1] ) );
  INV U2081 ( .IN(\mult_77/FS_1/TEMP_P[0][1][0] ), .OUT(m2549) );
  INV U2082 ( .IN(m2550), .OUT(\mult_77/FS_1/P[0][1][1] ) );
  INV U2083 ( .IN(\mult_76/FS_1/TEMP_P[0][1][0] ), .OUT(m2527) );
  INV U2084 ( .IN(m2528), .OUT(\mult_76/FS_1/P[0][1][1] ) );
  INV U2085 ( .IN(\mult_74/FS_1/TEMP_P[0][1][0] ), .OUT(m2506) );
  INV U2086 ( .IN(m2507), .OUT(\mult_74/FS_1/P[0][1][1] ) );
  INV U2087 ( .IN(\mult_72/FS_1/TEMP_P[0][1][0] ), .OUT(m2486) );
  INV U2088 ( .IN(m2487), .OUT(\mult_72/FS_1/P[0][1][1] ) );
  INV U2089 ( .IN(\mult_71/FS_1/TEMP_P[0][1][0] ), .OUT(m2464) );
  INV U2090 ( .IN(m2465), .OUT(\mult_71/FS_1/P[0][1][1] ) );
  INV U2091 ( .IN(m2595), .OUT(\mult_83/FS_1/P[0][1][3] ) );
  INV U2092 ( .IN(\mult_83/FS_1/P[0][1][3] ), .OUT(m2596) );
  INV U2093 ( .IN(m2597), .OUT(\mult_83/FS_1/TEMP_P[0][2][0] ) );
  INV U2094 ( .IN(\mult_83/FS_1/TEMP_P[0][2][0] ), .OUT(m2598) );
  INV U2095 ( .IN(m2599), .OUT(\mult_83/FS_1/P[0][2][1] ) );
  INV U2096 ( .IN(\mult_83/FS_1/P[0][2][1] ), .OUT(m2600) );
  INV U2097 ( .IN(\mult_83/FS_1/P[0][1][1] ), .OUT(m2592) );
  INV U2098 ( .IN(m2593), .OUT(\mult_83/FS_1/P[0][1][2] ) );
  INV U2099 ( .IN(\mult_83/FS_1/P[0][1][2] ), .OUT(m2594) );
  INV U2100 ( .IN(m2430), .OUT(\mult_82/FS_1/TEMP_P[0][2][0] ) );
  INV U2101 ( .IN(\mult_82/FS_1/TEMP_P[0][2][0] ), .OUT(m2431) );
  INV U2102 ( .IN(\mult_82/FS_1/P[0][1][1] ), .OUT(m2423) );
  INV U2103 ( .IN(m2424), .OUT(\mult_82/FS_1/P[0][1][2] ) );
  INV U2104 ( .IN(\mult_82/FS_1/P[0][1][2] ), .OUT(m2425) );
  INV U2105 ( .IN(m2578), .OUT(\mult_80/FS_1/TEMP_P[0][2][0] ) );
  INV U2106 ( .IN(\mult_80/FS_1/TEMP_P[0][2][0] ), .OUT(m2579) );
  INV U2107 ( .IN(\mult_80/FS_1/P[0][1][1] ), .OUT(m2571) );
  INV U2108 ( .IN(m2572), .OUT(\mult_80/FS_1/P[0][1][2] ) );
  INV U2109 ( .IN(\mult_80/FS_1/P[0][1][2] ), .OUT(m2573) );
  INV U2110 ( .IN(m2554), .OUT(\mult_77/FS_1/P[0][1][3] ) );
  INV U2111 ( .IN(\mult_77/FS_1/P[0][1][3] ), .OUT(m2555) );
  INV U2112 ( .IN(m2556), .OUT(\mult_77/FS_1/TEMP_P[0][2][0] ) );
  INV U2113 ( .IN(\mult_77/FS_1/TEMP_P[0][2][0] ), .OUT(m2557) );
  INV U2114 ( .IN(m2558), .OUT(\mult_77/FS_1/P[0][2][1] ) );
  INV U2115 ( .IN(\mult_77/FS_1/P[0][2][1] ), .OUT(m2559) );
  INV U2116 ( .IN(\mult_77/FS_1/P[0][1][1] ), .OUT(m2551) );
  INV U2117 ( .IN(m2552), .OUT(\mult_77/FS_1/P[0][1][2] ) );
  INV U2118 ( .IN(\mult_77/FS_1/P[0][1][2] ), .OUT(m2553) );
  INV U2119 ( .IN(m2536), .OUT(\mult_76/FS_1/TEMP_P[0][2][0] ) );
  INV U2120 ( .IN(\mult_76/FS_1/TEMP_P[0][2][0] ), .OUT(m2537) );
  INV U2121 ( .IN(\mult_76/FS_1/P[0][1][1] ), .OUT(m2529) );
  INV U2122 ( .IN(m2530), .OUT(\mult_76/FS_1/P[0][1][2] ) );
  INV U2123 ( .IN(\mult_76/FS_1/P[0][1][2] ), .OUT(m2531) );
  INV U2124 ( .IN(m2515), .OUT(\mult_74/FS_1/TEMP_P[0][2][0] ) );
  INV U2125 ( .IN(\mult_74/FS_1/TEMP_P[0][2][0] ), .OUT(m2516) );
  INV U2126 ( .IN(\mult_74/FS_1/P[0][1][1] ), .OUT(m2508) );
  INV U2127 ( .IN(m2509), .OUT(\mult_74/FS_1/P[0][1][2] ) );
  INV U2128 ( .IN(\mult_74/FS_1/P[0][1][2] ), .OUT(m2510) );
  INV U2129 ( .IN(m2491), .OUT(\mult_72/FS_1/P[0][1][3] ) );
  INV U2130 ( .IN(\mult_72/FS_1/P[0][1][3] ), .OUT(m2492) );
  INV U2131 ( .IN(m2493), .OUT(\mult_72/FS_1/TEMP_P[0][2][0] ) );
  INV U2132 ( .IN(\mult_72/FS_1/TEMP_P[0][2][0] ), .OUT(m2494) );
  INV U2133 ( .IN(m2495), .OUT(\mult_72/FS_1/P[0][2][1] ) );
  INV U2134 ( .IN(\mult_72/FS_1/P[0][2][1] ), .OUT(m2496) );
  INV U2135 ( .IN(\mult_72/FS_1/P[0][1][1] ), .OUT(m2488) );
  INV U2136 ( .IN(m2489), .OUT(\mult_72/FS_1/P[0][1][2] ) );
  INV U2137 ( .IN(\mult_72/FS_1/P[0][1][2] ), .OUT(m2490) );
  INV U2138 ( .IN(m2473), .OUT(\mult_71/FS_1/TEMP_P[0][2][0] ) );
  INV U2139 ( .IN(\mult_71/FS_1/TEMP_P[0][2][0] ), .OUT(m2474) );
  INV U2140 ( .IN(\mult_71/FS_1/P[0][1][1] ), .OUT(m2466) );
  INV U2141 ( .IN(m2467), .OUT(\mult_71/FS_1/P[0][1][2] ) );
  INV U2142 ( .IN(\mult_71/FS_1/P[0][1][2] ), .OUT(m2468) );
  INV U2143 ( .IN(\mult_69/FS_1/TEMP_P[0][0][0] ), .OUT(m2435) );
  INV U2144 ( .IN(m2436), .OUT(\mult_69/FS_1/P[0][0][1] ) );
  INV U2145 ( .IN(\mult_69/FS_1/P[0][0][1] ), .OUT(m2437) );
  INV U2146 ( .IN(m2438), .OUT(\mult_69/FS_1/P[0][0][2] ) );
  INV U2147 ( .IN(\mult_69/FS_1/P[0][0][2] ), .OUT(m2439) );
  INV U2148 ( .IN(m2440), .OUT(\mult_69/FS_1/P[0][0][3] ) );
  INV U2149 ( .IN(\mult_69/FS_1/P[0][0][3] ), .OUT(m2441) );
  INV U2150 ( .IN(m2442), .OUT(\mult_69/FS_1/TEMP_P[0][1][0] ) );
  INV U2151 ( .IN(\mult_69/FS_1/TEMP_P[0][1][0] ), .OUT(m2443) );
  INV U2152 ( .IN(m2444), .OUT(\mult_69/FS_1/P[0][1][1] ) );
  INV U2153 ( .IN(m2452), .OUT(\mult_69/FS_1/TEMP_P[0][2][0] ) );
  INV U2154 ( .IN(\mult_69/FS_1/TEMP_P[0][2][0] ), .OUT(m2453) );
  INV U2155 ( .IN(\mult_69/FS_1/P[0][1][1] ), .OUT(m2445) );
  INV U2156 ( .IN(m2446), .OUT(\mult_69/FS_1/P[0][1][2] ) );
  INV U2157 ( .IN(\mult_69/FS_1/P[0][1][2] ), .OUT(m2447) );
  INV U2158 ( .IN(\mult_82/A_not[7] ), .OUT(\mult_82/A1[8] ) );
  INV U2159 ( .IN(\mult_82/A_notx [6]), .OUT(\mult_82/A1[7] ) );
  INV U2160 ( .IN(\mult_82/A_notx [5]), .OUT(\mult_82/ab[5][3] ) );
  INV U2161 ( .IN(\mult_82/A_notx [4]), .OUT(\mult_82/ab[4][3] ) );
  INV U2162 ( .IN(\mult_82/A_notx [3]), .OUT(\mult_82/ab[3][3] ) );
  INV U2163 ( .IN(\mult_82/A_notx [2]), .OUT(\mult_82/ab[2][3] ) );
  INV U2164 ( .IN(\mult_82/A_notx [1]), .OUT(\mult_82/ab[1][3] ) );
  INV U2165 ( .IN(\mult_82/A_notx [0]), .OUT(\mult_82/ab[0][3] ) );
  INV U2166 ( .IN(\mult_82/A_notx [6]), .OUT(\mult_82/ab[6][0] ) );
  INV U2167 ( .IN(\mult_82/A_notx [5]), .OUT(\mult_82/ab[5][0] ) );
  INV U2168 ( .IN(\mult_82/A_notx [4]), .OUT(\mult_82/ab[4][0] ) );
  INV U2169 ( .IN(\mult_82/A_notx [3]), .OUT(\mult_82/ab[3][0] ) );
  INV U2170 ( .IN(\mult_82/A_notx [2]), .OUT(\mult_82/A1[0] ) );
  INV U2171 ( .IN(\mult_82/A_notx [1]), .OUT(N85) );
  INV U2172 ( .IN(\mult_82/A_notx [0]), .OUT(N84) );
  INV U2173 ( .IN(\mult_82/A_not[7] ), .OUT(\mult_82/ab[7][0] ) );
  INV U2174 ( .IN(\mult_69/A_not[7] ), .OUT(\mult_69/ab[7][2] ) );
  INV U2175 ( .IN(\mult_69/A_notx [6]), .OUT(\mult_69/ab[6][2] ) );
  INV U2176 ( .IN(\mult_69/A_notx [5]), .OUT(\mult_69/ab[5][2] ) );
  INV U2177 ( .IN(\mult_69/A_notx [4]), .OUT(\mult_69/ab[4][2] ) );
  INV U2178 ( .IN(\mult_69/A_notx [3]), .OUT(\mult_69/ab[3][2] ) );
  INV U2179 ( .IN(\mult_69/A_notx [2]), .OUT(\mult_69/ab[2][2] ) );
  INV U2180 ( .IN(\mult_69/A_notx [1]), .OUT(\mult_69/ab[1][2] ) );
  INV U2181 ( .IN(\mult_69/A_notx [0]), .OUT(\mult_69/ab[0][2] ) );
  INV U2182 ( .IN(\mult_69/A_notx [6]), .OUT(\mult_69/ab[6][1] ) );
  INV U2183 ( .IN(\mult_69/A_notx [5]), .OUT(\mult_69/ab[5][1] ) );
  INV U2184 ( .IN(\mult_69/A_notx [4]), .OUT(\mult_69/ab[4][1] ) );
  INV U2185 ( .IN(\mult_69/A_notx [3]), .OUT(\mult_69/ab[3][1] ) );
  INV U2186 ( .IN(\mult_69/A_notx [2]), .OUT(\mult_69/ab[2][1] ) );
  INV U2187 ( .IN(\mult_69/A_notx [1]), .OUT(\mult_69/ab[1][1] ) );
  INV U2188 ( .IN(\mult_69/A_notx [0]), .OUT(\mult_69/ab[0][1] ) );
  INV U2189 ( .IN(\mult_69/A_notx [6]), .OUT(\mult_69/ab[6][0] ) );
  INV U2190 ( .IN(\mult_69/A_notx [5]), .OUT(\mult_69/ab[5][0] ) );
  INV U2191 ( .IN(\mult_69/A_notx [4]), .OUT(\mult_69/ab[4][0] ) );
  INV U2192 ( .IN(\mult_69/A_notx [3]), .OUT(\mult_69/ab[3][0] ) );
  INV U2193 ( .IN(\mult_69/A_notx [2]), .OUT(\mult_69/ab[2][0] ) );
  INV U2194 ( .IN(\mult_69/A_notx [1]), .OUT(\mult_69/ab[1][0] ) );
  INV U2195 ( .IN(\mult_69/A_notx [0]), .OUT(N3) );
  INV U2196 ( .IN(\mult_69/A_not[7] ), .OUT(\mult_69/ab[7][0] ) );
  INV U2197 ( .IN(\mult_69/A_not[7] ), .OUT(\mult_69/ab[7][1] ) );
  INV U2198 ( .IN(\mult_71/A_not[7] ), .OUT(\mult_71/A1[8] ) );
  INV U2199 ( .IN(\mult_71/A_notx [6]), .OUT(\mult_71/A1[7] ) );
  INV U2200 ( .IN(\mult_71/A_notx [5]), .OUT(\mult_71/ab[5][3] ) );
  INV U2201 ( .IN(\mult_71/A_notx [4]), .OUT(\mult_71/ab[4][3] ) );
  INV U2202 ( .IN(\mult_71/A_notx [3]), .OUT(\mult_71/ab[3][3] ) );
  INV U2203 ( .IN(\mult_71/A_notx [2]), .OUT(\mult_71/ab[2][3] ) );
  INV U2204 ( .IN(\mult_71/A_notx [1]), .OUT(\mult_71/ab[1][3] ) );
  INV U2205 ( .IN(\mult_71/A_notx [0]), .OUT(\mult_71/ab[0][3] ) );
  INV U2206 ( .IN(\mult_71/A_notx [6]), .OUT(\mult_71/ab[6][0] ) );
  INV U2207 ( .IN(\mult_71/A_notx [5]), .OUT(\mult_71/ab[5][0] ) );
  INV U2208 ( .IN(\mult_71/A_notx [4]), .OUT(\mult_71/ab[4][0] ) );
  INV U2209 ( .IN(\mult_71/A_notx [3]), .OUT(\mult_71/ab[3][0] ) );
  INV U2210 ( .IN(\mult_71/A_notx [2]), .OUT(\mult_71/A1[0] ) );
  INV U2211 ( .IN(\mult_71/A_notx [1]), .OUT(N15) );
  INV U2212 ( .IN(\mult_71/A_notx [0]), .OUT(N14) );
  INV U2213 ( .IN(\mult_71/A_not[7] ), .OUT(\mult_71/ab[7][0] ) );
  INV U2214 ( .IN(\mult_72/A_not[7] ), .OUT(\mult_72/ab[7][3] ) );
  INV U2215 ( .IN(\mult_72/A_notx [6]), .OUT(\mult_72/ab[6][3] ) );
  INV U2216 ( .IN(\mult_72/A_notx [5]), .OUT(\mult_72/ab[5][3] ) );
  INV U2217 ( .IN(\mult_72/A_notx [4]), .OUT(\mult_72/ab[4][3] ) );
  INV U2218 ( .IN(\mult_72/A_notx [3]), .OUT(\mult_72/ab[3][3] ) );
  INV U2219 ( .IN(\mult_72/A_notx [2]), .OUT(\mult_72/ab[2][3] ) );
  INV U2220 ( .IN(\mult_72/A_notx [1]), .OUT(\mult_72/ab[1][3] ) );
  INV U2221 ( .IN(\mult_72/A_notx [0]), .OUT(\mult_72/ab[0][3] ) );
  INV U2222 ( .IN(\mult_72/A_notx [6]), .OUT(\mult_72/ab[6][2] ) );
  INV U2223 ( .IN(\mult_72/A_notx [5]), .OUT(\mult_72/ab[5][2] ) );
  INV U2224 ( .IN(\mult_72/A_notx [4]), .OUT(\mult_72/ab[4][2] ) );
  INV U2225 ( .IN(\mult_72/A_notx [3]), .OUT(\mult_72/ab[3][2] ) );
  INV U2226 ( .IN(\mult_72/A_notx [2]), .OUT(\mult_72/ab[2][2] ) );
  INV U2227 ( .IN(\mult_72/A_notx [1]), .OUT(\mult_72/ab[1][2] ) );
  INV U2228 ( .IN(\mult_72/A_notx [0]), .OUT(\mult_72/A1[0] ) );
  INV U2229 ( .IN(\mult_72/A_not[7] ), .OUT(\mult_72/ab[7][2] ) );
  INV U2230 ( .IN(\mult_74/A_not[7] ), .OUT(\mult_74/ab[7][2] ) );
  INV U2231 ( .IN(\mult_74/A_notx [6]), .OUT(\mult_74/ab[6][2] ) );
  INV U2232 ( .IN(\mult_74/A_notx [5]), .OUT(\mult_74/ab[5][2] ) );
  INV U2233 ( .IN(\mult_74/A_notx [4]), .OUT(\mult_74/ab[4][2] ) );
  INV U2234 ( .IN(\mult_74/A_notx [3]), .OUT(\mult_74/ab[3][2] ) );
  INV U2235 ( .IN(\mult_74/A_notx [2]), .OUT(\mult_74/ab[2][2] ) );
  INV U2236 ( .IN(\mult_74/A_notx [1]), .OUT(\mult_74/ab[1][2] ) );
  INV U2237 ( .IN(\mult_74/A_notx [0]), .OUT(\mult_74/ab[0][2] ) );
  INV U2238 ( .IN(\mult_74/A_notx [6]), .OUT(\mult_74/ab[6][1] ) );
  INV U2239 ( .IN(\mult_74/A_notx [5]), .OUT(\mult_74/ab[5][1] ) );
  INV U2240 ( .IN(\mult_74/A_notx [4]), .OUT(\mult_74/ab[4][1] ) );
  INV U2241 ( .IN(\mult_74/A_notx [3]), .OUT(\mult_74/ab[3][1] ) );
  INV U2242 ( .IN(\mult_74/A_notx [2]), .OUT(\mult_74/ab[2][1] ) );
  INV U2243 ( .IN(\mult_74/A_notx [1]), .OUT(\mult_74/ab[1][1] ) );
  INV U2244 ( .IN(\mult_74/A_notx [0]), .OUT(\mult_74/ab[0][1] ) );
  INV U2245 ( .IN(\mult_74/A_notx [6]), .OUT(\mult_74/ab[6][0] ) );
  INV U2246 ( .IN(\mult_74/A_notx [5]), .OUT(\mult_74/ab[5][0] ) );
  INV U2247 ( .IN(\mult_74/A_notx [4]), .OUT(\mult_74/ab[4][0] ) );
  INV U2248 ( .IN(\mult_74/A_notx [3]), .OUT(\mult_74/ab[3][0] ) );
  INV U2249 ( .IN(\mult_74/A_notx [2]), .OUT(\mult_74/ab[2][0] ) );
  INV U2250 ( .IN(\mult_74/A_notx [1]), .OUT(\mult_74/ab[1][0] ) );
  INV U2251 ( .IN(\mult_74/A_notx [0]), .OUT(N38) );
  INV U2252 ( .IN(\mult_74/A_not[7] ), .OUT(\mult_74/ab[7][0] ) );
  INV U2253 ( .IN(\mult_74/A_not[7] ), .OUT(\mult_74/ab[7][1] ) );
  INV U2254 ( .IN(\mult_76/A_not[7] ), .OUT(\mult_76/A1[8] ) );
  INV U2255 ( .IN(\mult_76/A_notx [6]), .OUT(\mult_76/A1[7] ) );
  INV U2256 ( .IN(\mult_76/A_notx [5]), .OUT(\mult_76/ab[5][3] ) );
  INV U2257 ( .IN(\mult_76/A_notx [4]), .OUT(\mult_76/ab[4][3] ) );
  INV U2258 ( .IN(\mult_76/A_notx [3]), .OUT(\mult_76/ab[3][3] ) );
  INV U2259 ( .IN(\mult_76/A_notx [2]), .OUT(\mult_76/ab[2][3] ) );
  INV U2260 ( .IN(\mult_76/A_notx [1]), .OUT(\mult_76/ab[1][3] ) );
  INV U2261 ( .IN(\mult_76/A_notx [0]), .OUT(\mult_76/ab[0][3] ) );
  INV U2262 ( .IN(\mult_76/A_notx [6]), .OUT(\mult_76/ab[6][0] ) );
  INV U2263 ( .IN(\mult_76/A_notx [5]), .OUT(\mult_76/ab[5][0] ) );
  INV U2264 ( .IN(\mult_76/A_notx [4]), .OUT(\mult_76/ab[4][0] ) );
  INV U2265 ( .IN(\mult_76/A_notx [3]), .OUT(\mult_76/ab[3][0] ) );
  INV U2266 ( .IN(\mult_76/A_notx [2]), .OUT(\mult_76/A1[0] ) );
  INV U2267 ( .IN(\mult_76/A_notx [1]), .OUT(N50) );
  INV U2268 ( .IN(\mult_76/A_notx [0]), .OUT(N49) );
  INV U2269 ( .IN(\mult_76/A_not[7] ), .OUT(\mult_76/ab[7][0] ) );
  INV U2270 ( .IN(\mult_77/A_not[7] ), .OUT(\mult_77/ab[7][3] ) );
  INV U2271 ( .IN(\mult_77/A_notx [6]), .OUT(\mult_77/ab[6][3] ) );
  INV U2272 ( .IN(\mult_77/A_notx [5]), .OUT(\mult_77/ab[5][3] ) );
  INV U2273 ( .IN(\mult_77/A_notx [4]), .OUT(\mult_77/ab[4][3] ) );
  INV U2274 ( .IN(\mult_77/A_notx [3]), .OUT(\mult_77/ab[3][3] ) );
  INV U2275 ( .IN(\mult_77/A_notx [2]), .OUT(\mult_77/ab[2][3] ) );
  INV U2276 ( .IN(\mult_77/A_notx [1]), .OUT(\mult_77/ab[1][3] ) );
  INV U2277 ( .IN(\mult_77/A_notx [0]), .OUT(\mult_77/ab[0][3] ) );
  INV U2278 ( .IN(\mult_77/A_notx [6]), .OUT(\mult_77/ab[6][2] ) );
  INV U2279 ( .IN(\mult_77/A_notx [5]), .OUT(\mult_77/ab[5][2] ) );
  INV U2280 ( .IN(\mult_77/A_notx [4]), .OUT(\mult_77/ab[4][2] ) );
  INV U2281 ( .IN(\mult_77/A_notx [3]), .OUT(\mult_77/ab[3][2] ) );
  INV U2282 ( .IN(\mult_77/A_notx [2]), .OUT(\mult_77/ab[2][2] ) );
  INV U2283 ( .IN(\mult_77/A_notx [1]), .OUT(\mult_77/ab[1][2] ) );
  INV U2284 ( .IN(\mult_77/A_notx [0]), .OUT(\mult_77/A1[0] ) );
  INV U2285 ( .IN(\mult_77/A_not[7] ), .OUT(\mult_77/ab[7][2] ) );
  INV U2286 ( .IN(\mult_80/A_not[7] ), .OUT(\mult_80/ab[7][2] ) );
  INV U2287 ( .IN(\mult_80/A_notx [6]), .OUT(\mult_80/ab[6][2] ) );
  INV U2288 ( .IN(\mult_80/A_notx [5]), .OUT(\mult_80/ab[5][2] ) );
  INV U2289 ( .IN(\mult_80/A_notx [4]), .OUT(\mult_80/ab[4][2] ) );
  INV U2290 ( .IN(\mult_80/A_notx [3]), .OUT(\mult_80/ab[3][2] ) );
  INV U2291 ( .IN(\mult_80/A_notx [2]), .OUT(\mult_80/ab[2][2] ) );
  INV U2292 ( .IN(\mult_80/A_notx [1]), .OUT(\mult_80/ab[1][2] ) );
  INV U2293 ( .IN(\mult_80/A_notx [0]), .OUT(\mult_80/ab[0][2] ) );
  INV U2294 ( .IN(\mult_80/A_notx [6]), .OUT(\mult_80/ab[6][1] ) );
  INV U2295 ( .IN(\mult_80/A_notx [5]), .OUT(\mult_80/ab[5][1] ) );
  INV U2296 ( .IN(\mult_80/A_notx [4]), .OUT(\mult_80/ab[4][1] ) );
  INV U2297 ( .IN(\mult_80/A_notx [3]), .OUT(\mult_80/ab[3][1] ) );
  INV U2298 ( .IN(\mult_80/A_notx [2]), .OUT(\mult_80/ab[2][1] ) );
  INV U2299 ( .IN(\mult_80/A_notx [1]), .OUT(\mult_80/ab[1][1] ) );
  INV U2300 ( .IN(\mult_80/A_notx [0]), .OUT(\mult_80/ab[0][1] ) );
  INV U2301 ( .IN(\mult_80/A_notx [6]), .OUT(\mult_80/ab[6][0] ) );
  INV U2302 ( .IN(\mult_80/A_notx [5]), .OUT(\mult_80/ab[5][0] ) );
  INV U2303 ( .IN(\mult_80/A_notx [4]), .OUT(\mult_80/ab[4][0] ) );
  INV U2304 ( .IN(\mult_80/A_notx [3]), .OUT(\mult_80/ab[3][0] ) );
  INV U2305 ( .IN(\mult_80/A_notx [2]), .OUT(\mult_80/ab[2][0] ) );
  INV U2306 ( .IN(\mult_80/A_notx [1]), .OUT(\mult_80/ab[1][0] ) );
  INV U2307 ( .IN(\mult_80/A_notx [0]), .OUT(N73) );
  INV U2308 ( .IN(\mult_80/A_not[7] ), .OUT(\mult_80/ab[7][0] ) );
  INV U2309 ( .IN(\mult_80/A_not[7] ), .OUT(\mult_80/ab[7][1] ) );
  INV U2310 ( .IN(\mult_83/A_not[7] ), .OUT(\mult_83/ab[7][3] ) );
  INV U2311 ( .IN(\mult_83/A_notx [6]), .OUT(\mult_83/ab[6][3] ) );
  INV U2312 ( .IN(\mult_83/A_notx [5]), .OUT(\mult_83/ab[5][3] ) );
  INV U2313 ( .IN(\mult_83/A_notx [4]), .OUT(\mult_83/ab[4][3] ) );
  INV U2314 ( .IN(\mult_83/A_notx [3]), .OUT(\mult_83/ab[3][3] ) );
  INV U2315 ( .IN(\mult_83/A_notx [2]), .OUT(\mult_83/ab[2][3] ) );
  INV U2316 ( .IN(\mult_83/A_notx [1]), .OUT(\mult_83/ab[1][3] ) );
  INV U2317 ( .IN(\mult_83/A_notx [0]), .OUT(\mult_83/ab[0][3] ) );
  INV U2318 ( .IN(\mult_83/A_notx [6]), .OUT(\mult_83/ab[6][2] ) );
  INV U2319 ( .IN(\mult_83/A_notx [5]), .OUT(\mult_83/ab[5][2] ) );
  INV U2320 ( .IN(\mult_83/A_notx [4]), .OUT(\mult_83/ab[4][2] ) );
  INV U2321 ( .IN(\mult_83/A_notx [3]), .OUT(\mult_83/ab[3][2] ) );
  INV U2322 ( .IN(\mult_83/A_notx [2]), .OUT(\mult_83/ab[2][2] ) );
  INV U2323 ( .IN(\mult_83/A_notx [1]), .OUT(\mult_83/ab[1][2] ) );
  INV U2324 ( .IN(\mult_83/A_notx [0]), .OUT(\mult_83/A1[0] ) );
  INV U2325 ( .IN(\mult_83/A_not[7] ), .OUT(\mult_83/ab[7][2] ) );
  INV U2326 ( .IN(\mult_82/FS_1/G[1][0][1] ), .OUT(m2433) );
  INV U2327 ( .IN(\mult_80/FS_1/G[1][0][1] ), .OUT(m2580) );
  INV U2328 ( .IN(\mult_76/FS_1/G[1][0][1] ), .OUT(m2539) );
  INV U2329 ( .IN(\mult_74/FS_1/G[1][0][1] ), .OUT(m2517) );
  INV U2330 ( .IN(\mult_71/FS_1/G[1][0][1] ), .OUT(m2476) );
  NAND2 U2331 ( .A(\mult_82/FS_1/C[1][2][0] ), .B(
        \mult_82/FS_1/TEMP_P[0][2][0] ), .OUT(m2432) );
  INV U2332 ( .IN(\mult_82/FS_1/G[0][1][3] ), .OUT(m2429) );
  INV U2333 ( .IN(\mult_80/FS_1/G[0][1][3] ), .OUT(m2577) );
  NAND2 U2334 ( .A(\mult_76/FS_1/C[1][2][0] ), .B(
        \mult_76/FS_1/TEMP_P[0][2][0] ), .OUT(m2538) );
  INV U2335 ( .IN(\mult_76/FS_1/G[0][1][3] ), .OUT(m2535) );
  INV U2336 ( .IN(\mult_74/FS_1/G[0][1][3] ), .OUT(m2514) );
  NAND2 U2337 ( .A(\mult_71/FS_1/C[1][2][0] ), .B(
        \mult_71/FS_1/TEMP_P[0][2][0] ), .OUT(m2475) );
  INV U2338 ( .IN(\mult_71/FS_1/G[0][1][3] ), .OUT(m2472) );
  INV U2339 ( .IN(\mult_69/FS_1/G[1][0][1] ), .OUT(m2454) );
  INV U2340 ( .IN(\mult_69/FS_1/G[0][1][3] ), .OUT(m2451) );
  NOR2 U2341 ( .A(m1316), .B(m1317), .OUT(\mult_82/A2[7] ) );
  NOR2 U2342 ( .A(m1318), .B(m1319), .OUT(\mult_69/A2[8] ) );
  NOR2 U2343 ( .A(m1320), .B(m1321), .OUT(\mult_69/A2[7] ) );
  NOR2 U2344 ( .A(m1322), .B(m1323), .OUT(\mult_71/A2[7] ) );
  NOR2 U2345 ( .A(m1324), .B(m1325), .OUT(\mult_72/A2[9] ) );
  NOR2 U2346 ( .A(m1326), .B(m1327), .OUT(\mult_74/A2[8] ) );
  NOR2 U2347 ( .A(m1328), .B(m1329), .OUT(\mult_74/A2[7] ) );
  NOR2 U2348 ( .A(m1330), .B(m1331), .OUT(\mult_76/A2[7] ) );
  NOR2 U2349 ( .A(m1332), .B(m1333), .OUT(\mult_77/A2[9] ) );
  NOR2 U2350 ( .A(m1334), .B(m1335), .OUT(\mult_80/A2[8] ) );
  NOR2 U2351 ( .A(m1336), .B(m1337), .OUT(\mult_80/A2[7] ) );
  NOR2 U2352 ( .A(m1338), .B(m1339), .OUT(\mult_83/A2[9] ) );
  OAI22 U2353 ( .A(m1340), .B(m1341), .C(m1342), .D(m1343), .OUT(N119) );
  NOR2 U2354 ( .A(\mult_83/ab[1][3] ), .B(\mult_83/ab[2][2] ), .OUT(m1344) );
  NOR2 U2355 ( .A(\mult_83/ab[2][3] ), .B(\mult_83/ab[3][2] ), .OUT(m1345) );
  NOR2 U2356 ( .A(\mult_83/ab[3][3] ), .B(\mult_83/ab[4][2] ), .OUT(m1346) );
  NOR2 U2357 ( .A(\mult_83/ab[4][3] ), .B(\mult_83/ab[5][2] ), .OUT(m1347) );
  NOR2 U2358 ( .A(\mult_83/ab[5][3] ), .B(\mult_83/ab[6][2] ), .OUT(m1348) );
  NOR2 U2359 ( .A(\mult_83/ab[6][3] ), .B(\mult_83/ab[7][2] ), .OUT(m1349) );
  NOR2 U2360 ( .A(\mult_82/ab[4][0] ), .B(m1351), .OUT(m1350) );
  NAND2 U2361 ( .A(m1353), .B(m1354), .OUT(m1352) );
  NAND2 U2362 ( .A(m1356), .B(m1357), .OUT(m1355) );
  NAND2 U2363 ( .A(m1359), .B(m1360), .OUT(m1358) );
  NOR2 U2364 ( .A(\mult_80/ab[1][2] ), .B(\mult_80/ab[2][1] ), .OUT(m1361) );
  NOR2 U2365 ( .A(\mult_80/ab[2][2] ), .B(\mult_80/ab[3][1] ), .OUT(m1362) );
  NOR2 U2366 ( .A(\mult_80/ab[3][2] ), .B(\mult_80/ab[4][1] ), .OUT(m1363) );
  NOR2 U2367 ( .A(\mult_80/ab[4][2] ), .B(\mult_80/ab[5][1] ), .OUT(m1364) );
  NOR2 U2368 ( .A(\mult_80/ab[5][2] ), .B(\mult_80/ab[6][1] ), .OUT(m1365) );
  NOR2 U2369 ( .A(\mult_80/ab[6][2] ), .B(\mult_80/ab[7][1] ), .OUT(m1366) );
  NAND2 U2370 ( .A(m1368), .B(m1369), .OUT(m1367) );
  NOR2 U2371 ( .A(\mult_80/ab[3][0] ), .B(m1371), .OUT(m1370) );
  NOR2 U2372 ( .A(\mult_80/ab[4][0] ), .B(m1373), .OUT(m1372) );
  NOR2 U2373 ( .A(\mult_80/ab[5][0] ), .B(m1375), .OUT(m1374) );
  NOR2 U2374 ( .A(\mult_80/ab[6][0] ), .B(m1377), .OUT(m1376) );
  NOR2 U2375 ( .A(\mult_80/ab[7][0] ), .B(m1379), .OUT(m1378) );
  NOR2 U2376 ( .A(\mult_77/ab[1][3] ), .B(\mult_77/ab[2][2] ), .OUT(m1380) );
  NOR2 U2377 ( .A(\mult_77/ab[2][3] ), .B(\mult_77/ab[3][2] ), .OUT(m1381) );
  NOR2 U2378 ( .A(\mult_77/ab[3][3] ), .B(\mult_77/ab[4][2] ), .OUT(m1382) );
  NOR2 U2379 ( .A(\mult_77/ab[4][3] ), .B(\mult_77/ab[5][2] ), .OUT(m1383) );
  NOR2 U2380 ( .A(\mult_77/ab[5][3] ), .B(\mult_77/ab[6][2] ), .OUT(m1384) );
  NOR2 U2381 ( .A(\mult_77/ab[6][3] ), .B(\mult_77/ab[7][2] ), .OUT(m1385) );
  NOR2 U2382 ( .A(\mult_76/ab[4][0] ), .B(m1387), .OUT(m1386) );
  NAND2 U2383 ( .A(m1389), .B(m1390), .OUT(m1388) );
  NAND2 U2384 ( .A(m1392), .B(m1393), .OUT(m1391) );
  NAND2 U2385 ( .A(m1395), .B(m1396), .OUT(m1394) );
  NOR2 U2386 ( .A(\mult_74/ab[1][2] ), .B(\mult_74/ab[2][1] ), .OUT(m1397) );
  NOR2 U2387 ( .A(\mult_74/ab[2][2] ), .B(\mult_74/ab[3][1] ), .OUT(m1398) );
  NOR2 U2388 ( .A(\mult_74/ab[3][2] ), .B(\mult_74/ab[4][1] ), .OUT(m1399) );
  NOR2 U2389 ( .A(\mult_74/ab[4][2] ), .B(\mult_74/ab[5][1] ), .OUT(m1400) );
  NOR2 U2390 ( .A(\mult_74/ab[5][2] ), .B(\mult_74/ab[6][1] ), .OUT(m1401) );
  NOR2 U2391 ( .A(\mult_74/ab[6][2] ), .B(\mult_74/ab[7][1] ), .OUT(m1402) );
  NAND2 U2392 ( .A(m1404), .B(m1405), .OUT(m1403) );
  NOR2 U2393 ( .A(\mult_74/ab[3][0] ), .B(m1407), .OUT(m1406) );
  NOR2 U2394 ( .A(\mult_74/ab[4][0] ), .B(m1409), .OUT(m1408) );
  NOR2 U2395 ( .A(\mult_74/ab[5][0] ), .B(m1411), .OUT(m1410) );
  NOR2 U2396 ( .A(\mult_74/ab[6][0] ), .B(m1413), .OUT(m1412) );
  NOR2 U2397 ( .A(\mult_74/ab[7][0] ), .B(m1415), .OUT(m1414) );
  NOR2 U2398 ( .A(\mult_72/ab[1][3] ), .B(\mult_72/ab[2][2] ), .OUT(m1416) );
  NOR2 U2399 ( .A(\mult_72/ab[2][3] ), .B(\mult_72/ab[3][2] ), .OUT(m1417) );
  NOR2 U2400 ( .A(\mult_72/ab[3][3] ), .B(\mult_72/ab[4][2] ), .OUT(m1418) );
  NOR2 U2401 ( .A(\mult_72/ab[4][3] ), .B(\mult_72/ab[5][2] ), .OUT(m1419) );
  NOR2 U2402 ( .A(\mult_72/ab[5][3] ), .B(\mult_72/ab[6][2] ), .OUT(m1420) );
  NOR2 U2403 ( .A(\mult_72/ab[6][3] ), .B(\mult_72/ab[7][2] ), .OUT(m1421) );
  NOR2 U2404 ( .A(\mult_71/ab[4][0] ), .B(m1423), .OUT(m1422) );
  NAND2 U2405 ( .A(m1425), .B(m1426), .OUT(m1424) );
  NAND2 U2406 ( .A(m1428), .B(m1429), .OUT(m1427) );
  NAND2 U2407 ( .A(m1431), .B(m1432), .OUT(m1430) );
  NOR2 U2408 ( .A(\mult_69/ab[1][2] ), .B(\mult_69/ab[2][1] ), .OUT(m1433) );
  NOR2 U2409 ( .A(\mult_69/ab[2][2] ), .B(\mult_69/ab[3][1] ), .OUT(m1434) );
  NOR2 U2410 ( .A(\mult_69/ab[3][2] ), .B(\mult_69/ab[4][1] ), .OUT(m1435) );
  NOR2 U2411 ( .A(\mult_69/ab[4][2] ), .B(\mult_69/ab[5][1] ), .OUT(m1436) );
  NOR2 U2412 ( .A(\mult_69/ab[5][2] ), .B(\mult_69/ab[6][1] ), .OUT(m1437) );
  NOR2 U2413 ( .A(\mult_69/ab[6][2] ), .B(\mult_69/ab[7][1] ), .OUT(m1438) );
  NAND2 U2414 ( .A(m1440), .B(m1441), .OUT(m1439) );
  NOR2 U2415 ( .A(\mult_69/ab[3][0] ), .B(m1443), .OUT(m1442) );
  NOR2 U2416 ( .A(\mult_69/ab[4][0] ), .B(m1445), .OUT(m1444) );
  NOR2 U2417 ( .A(\mult_69/ab[5][0] ), .B(m1447), .OUT(m1446) );
  NOR2 U2418 ( .A(\mult_69/ab[6][0] ), .B(m1449), .OUT(m1448) );
  NOR2 U2419 ( .A(\mult_69/ab[7][0] ), .B(m1451), .OUT(m1450) );
  NOR2 U2420 ( .A(\PR_mul[14][3] ), .B(\PR_add[12][3] ), .OUT(m1452) );
  NOR2 U2421 ( .A(\PR_mul[14][4] ), .B(\PR_add[12][4] ), .OUT(m1453) );
  NOR2 U2422 ( .A(\PR_mul[14][5] ), .B(\PR_add[12][5] ), .OUT(m1454) );
  NOR2 U2423 ( .A(\PR_mul[14][6] ), .B(\PR_add[12][6] ), .OUT(m1455) );
  NOR2 U2424 ( .A(\PR_mul[14][7] ), .B(\PR_add[12][7] ), .OUT(m1456) );
  NOR2 U2425 ( .A(\PR_mul[14][8] ), .B(\PR_add[12][8] ), .OUT(m1457) );
  NOR2 U2426 ( .A(\PR_mul[14][9] ), .B(\PR_add[12][9] ), .OUT(m1458) );
  NOR2 U2427 ( .A(m1460), .B(m1461), .OUT(m1459) );
  NAND2 U2428 ( .A(\PR_add[12][16] ), .B(m1463), .OUT(m1462) );
  NAND2 U2429 ( .A(\PR_add[12][14] ), .B(m1465), .OUT(m1464) );
  NOR2 U2430 ( .A(m1467), .B(m1468), .OUT(m1466) );
  NAND2 U2431 ( .A(m1470), .B(\PR_add[12][10] ), .OUT(m1469) );
  NOR2 U2432 ( .A(\PR_mul[13][3] ), .B(\PR_add[11][3] ), .OUT(m1471) );
  NOR2 U2433 ( .A(\PR_mul[13][4] ), .B(\PR_add[11][4] ), .OUT(m1472) );
  NOR2 U2434 ( .A(\PR_mul[13][5] ), .B(\PR_add[11][5] ), .OUT(m1473) );
  NOR2 U2435 ( .A(\PR_mul[13][6] ), .B(\PR_add[11][6] ), .OUT(m1474) );
  NOR2 U2436 ( .A(\PR_mul[13][7] ), .B(\PR_add[11][7] ), .OUT(m1475) );
  NOR2 U2437 ( .A(\PR_mul[13][8] ), .B(\PR_add[11][8] ), .OUT(m1476) );
  NOR2 U2438 ( .A(\PR_mul[13][9] ), .B(\PR_add[11][9] ), .OUT(m1477) );
  NOR2 U2439 ( .A(\PR_mul[13][10] ), .B(\PR_add[11][10] ), .OUT(m1478) );
  NOR2 U2440 ( .A(\PR_mul[13][11] ), .B(\PR_add[11][11] ), .OUT(m1479) );
  NOR2 U2441 ( .A(m1481), .B(m1482), .OUT(m1480) );
  NAND2 U2442 ( .A(\PR_add[11][16] ), .B(m1484), .OUT(m1483) );
  NAND2 U2443 ( .A(m1486), .B(\PR_add[11][12] ), .OUT(m1485) );
  NOR2 U2444 ( .A(\PR_mul[12][1] ), .B(\PR_add[10][1] ), .OUT(m1487) );
  NOR2 U2445 ( .A(\PR_mul[12][2] ), .B(\PR_add[10][2] ), .OUT(m1488) );
  NOR2 U2446 ( .A(\PR_mul[12][3] ), .B(\PR_add[10][3] ), .OUT(m1489) );
  NOR2 U2447 ( .A(\PR_mul[12][4] ), .B(\PR_add[10][4] ), .OUT(m1490) );
  NOR2 U2448 ( .A(\PR_mul[12][5] ), .B(\PR_add[10][5] ), .OUT(m1491) );
  NOR2 U2449 ( .A(\PR_mul[12][6] ), .B(\PR_add[10][6] ), .OUT(m1492) );
  NOR2 U2450 ( .A(\PR_mul[12][7] ), .B(\PR_add[10][7] ), .OUT(m1493) );
  NOR2 U2451 ( .A(\PR_mul[12][8] ), .B(\PR_add[10][8] ), .OUT(m1494) );
  NOR2 U2452 ( .A(\PR_mul[12][9] ), .B(\PR_add[10][9] ), .OUT(m1495) );
  NOR2 U2453 ( .A(\PR_mul[12][10] ), .B(\PR_add[10][10] ), .OUT(m1496) );
  NOR2 U2454 ( .A(\PR_mul[12][11] ), .B(\PR_add[10][11] ), .OUT(m1497) );
  NOR2 U2455 ( .A(m1499), .B(m1500), .OUT(m1498) );
  NAND2 U2456 ( .A(\PR_add[10][16] ), .B(m1502), .OUT(m1501) );
  NAND2 U2457 ( .A(m1504), .B(\PR_add[10][12] ), .OUT(m1503) );
  NOR2 U2458 ( .A(\PR_mul[11][4] ), .B(\PR_add[9][4] ), .OUT(m1505) );
  NOR2 U2459 ( .A(\PR_mul[11][5] ), .B(\PR_add[9][5] ), .OUT(m1506) );
  NOR2 U2460 ( .A(\PR_mul[11][6] ), .B(\PR_add[9][6] ), .OUT(m1507) );
  NOR2 U2461 ( .A(\PR_mul[11][7] ), .B(\PR_add[9][7] ), .OUT(m1508) );
  NOR2 U2462 ( .A(\PR_mul[11][8] ), .B(\PR_add[9][8] ), .OUT(m1509) );
  NOR2 U2463 ( .A(\PR_mul[11][9] ), .B(\PR_add[9][9] ), .OUT(m1510) );
  NOR2 U2464 ( .A(\PR_mul[11][10] ), .B(\PR_add[9][10] ), .OUT(m1511) );
  NAND2 U2465 ( .A(m1513), .B(\PR_add[9][18] ), .OUT(m1512) );
  NAND2 U2466 ( .A(\PR_add[9][15] ), .B(m1515), .OUT(m1514) );
  NOR2 U2467 ( .A(m1517), .B(m1518), .OUT(m1516) );
  NAND2 U2468 ( .A(m1520), .B(\PR_add[9][11] ), .OUT(m1519) );
  NOR2 U2469 ( .A(\PR_mul[10][1] ), .B(\PR_add[8][1] ), .OUT(m1521) );
  NOR2 U2470 ( .A(\PR_mul[10][2] ), .B(\PR_add[8][2] ), .OUT(m1522) );
  NOR2 U2471 ( .A(\PR_mul[10][3] ), .B(\PR_add[8][3] ), .OUT(m1523) );
  NOR2 U2472 ( .A(\PR_mul[10][4] ), .B(\PR_add[8][4] ), .OUT(m1524) );
  NOR2 U2473 ( .A(\PR_mul[10][5] ), .B(\PR_add[8][5] ), .OUT(m1525) );
  NOR2 U2474 ( .A(\PR_mul[10][6] ), .B(\PR_add[8][6] ), .OUT(m1526) );
  NOR2 U2475 ( .A(\PR_mul[10][7] ), .B(\PR_add[8][7] ), .OUT(m1527) );
  NOR2 U2476 ( .A(\PR_mul[10][8] ), .B(\PR_add[8][8] ), .OUT(m1528) );
  NOR2 U2477 ( .A(\PR_mul[10][9] ), .B(\PR_add[8][9] ), .OUT(m1529) );
  NOR2 U2478 ( .A(\PR_mul[10][10] ), .B(\PR_add[8][10] ), .OUT(m1530) );
  NAND2 U2479 ( .A(m1532), .B(\PR_add[8][18] ), .OUT(m1531) );
  NAND2 U2480 ( .A(\PR_add[8][15] ), .B(m1534), .OUT(m1533) );
  NOR2 U2481 ( .A(m1536), .B(m1537), .OUT(m1535) );
  NAND2 U2482 ( .A(m1539), .B(\PR_add[8][11] ), .OUT(m1538) );
  NOR2 U2483 ( .A(\PR_mul[9][3] ), .B(\PR_add[7][3] ), .OUT(m1540) );
  NOR2 U2484 ( .A(\PR_mul[9][4] ), .B(\PR_add[7][4] ), .OUT(m1541) );
  NOR2 U2485 ( .A(\PR_mul[9][5] ), .B(\PR_add[7][5] ), .OUT(m1542) );
  NOR2 U2486 ( .A(\PR_mul[9][6] ), .B(\PR_add[7][6] ), .OUT(m1543) );
  NOR2 U2487 ( .A(\PR_mul[9][7] ), .B(\PR_add[7][7] ), .OUT(m1544) );
  NOR2 U2488 ( .A(\PR_mul[9][8] ), .B(\PR_add[7][8] ), .OUT(m1545) );
  NOR2 U2489 ( .A(\PR_mul[9][9] ), .B(\PR_add[7][9] ), .OUT(m1546) );
  NOR2 U2490 ( .A(m1548), .B(m1549), .OUT(m1547) );
  NAND2 U2491 ( .A(\PR_add[7][16] ), .B(m1551), .OUT(m1550) );
  NAND2 U2492 ( .A(\PR_add[7][14] ), .B(m1553), .OUT(m1552) );
  NOR2 U2493 ( .A(m1555), .B(m1556), .OUT(m1554) );
  NAND2 U2494 ( .A(m1558), .B(\PR_add[7][10] ), .OUT(m1557) );
  NOR2 U2495 ( .A(\PR_mul[8][3] ), .B(\PR_add[6][3] ), .OUT(m1559) );
  NOR2 U2496 ( .A(\PR_mul[8][4] ), .B(\PR_add[6][4] ), .OUT(m1560) );
  NOR2 U2497 ( .A(\PR_mul[8][5] ), .B(\PR_add[6][5] ), .OUT(m1561) );
  NOR2 U2498 ( .A(\PR_mul[8][6] ), .B(\PR_add[6][6] ), .OUT(m1562) );
  NOR2 U2499 ( .A(\PR_mul[8][7] ), .B(\PR_add[6][7] ), .OUT(m1563) );
  NOR2 U2500 ( .A(\PR_mul[8][8] ), .B(\PR_add[6][8] ), .OUT(m1564) );
  NOR2 U2501 ( .A(\PR_mul[8][9] ), .B(\PR_add[6][9] ), .OUT(m1565) );
  NOR2 U2502 ( .A(\PR_mul[8][10] ), .B(\PR_add[6][10] ), .OUT(m1566) );
  NOR2 U2503 ( .A(\PR_mul[8][11] ), .B(\PR_add[6][11] ), .OUT(m1567) );
  NOR2 U2504 ( .A(m1569), .B(m1570), .OUT(m1568) );
  NAND2 U2505 ( .A(\PR_add[6][16] ), .B(m1572), .OUT(m1571) );
  NAND2 U2506 ( .A(m1574), .B(\PR_add[6][12] ), .OUT(m1573) );
  NOR2 U2507 ( .A(\PR_mul[7][1] ), .B(\PR_add[5][1] ), .OUT(m1575) );
  NOR2 U2508 ( .A(\PR_mul[7][2] ), .B(\PR_add[5][2] ), .OUT(m1576) );
  NOR2 U2509 ( .A(\PR_mul[7][3] ), .B(\PR_add[5][3] ), .OUT(m1577) );
  NOR2 U2510 ( .A(\PR_mul[7][4] ), .B(\PR_add[5][4] ), .OUT(m1578) );
  NOR2 U2511 ( .A(\PR_mul[7][5] ), .B(\PR_add[5][5] ), .OUT(m1579) );
  NOR2 U2512 ( .A(\PR_mul[7][6] ), .B(\PR_add[5][6] ), .OUT(m1580) );
  NOR2 U2513 ( .A(\PR_mul[7][7] ), .B(\PR_add[5][7] ), .OUT(m1581) );
  NOR2 U2514 ( .A(\PR_mul[7][8] ), .B(\PR_add[5][8] ), .OUT(m1582) );
  NOR2 U2515 ( .A(\PR_mul[7][9] ), .B(\PR_add[5][9] ), .OUT(m1583) );
  NOR2 U2516 ( .A(\PR_mul[7][10] ), .B(\PR_add[5][10] ), .OUT(m1584) );
  NOR2 U2517 ( .A(\PR_mul[7][11] ), .B(\PR_add[5][11] ), .OUT(m1585) );
  NOR2 U2518 ( .A(m1587), .B(m1588), .OUT(m1586) );
  NAND2 U2519 ( .A(\PR_add[5][16] ), .B(m1590), .OUT(m1589) );
  NAND2 U2520 ( .A(m1592), .B(\PR_add[5][12] ), .OUT(m1591) );
  NOR2 U2521 ( .A(\PR_mul[6][4] ), .B(\PR_add[4][4] ), .OUT(m1593) );
  NOR2 U2522 ( .A(\PR_mul[6][5] ), .B(\PR_add[4][5] ), .OUT(m1594) );
  NOR2 U2523 ( .A(\PR_mul[6][6] ), .B(\PR_add[4][6] ), .OUT(m1595) );
  NOR2 U2524 ( .A(\PR_mul[6][7] ), .B(\PR_add[4][7] ), .OUT(m1596) );
  NOR2 U2525 ( .A(\PR_mul[6][8] ), .B(\PR_add[4][8] ), .OUT(m1597) );
  NOR2 U2526 ( .A(\PR_mul[6][9] ), .B(\PR_add[4][9] ), .OUT(m1598) );
  NOR2 U2527 ( .A(\PR_mul[6][10] ), .B(\PR_add[4][10] ), .OUT(m1599) );
  NAND2 U2528 ( .A(m1601), .B(\PR_add[4][18] ), .OUT(m1600) );
  NAND2 U2529 ( .A(\PR_add[4][15] ), .B(m1603), .OUT(m1602) );
  NOR2 U2530 ( .A(m1605), .B(m1606), .OUT(m1604) );
  NAND2 U2531 ( .A(m1608), .B(\PR_add[4][11] ), .OUT(m1607) );
  NOR2 U2532 ( .A(\PR_mul[5][1] ), .B(\PR_add[3][1] ), .OUT(m1609) );
  NOR2 U2533 ( .A(\PR_mul[5][2] ), .B(\PR_add[3][2] ), .OUT(m1610) );
  NOR2 U2534 ( .A(\PR_mul[5][3] ), .B(\PR_add[3][3] ), .OUT(m1611) );
  NOR2 U2535 ( .A(\PR_mul[5][4] ), .B(\PR_add[3][4] ), .OUT(m1612) );
  NOR2 U2536 ( .A(\PR_mul[5][5] ), .B(\PR_add[3][5] ), .OUT(m1613) );
  NOR2 U2537 ( .A(\PR_mul[5][6] ), .B(\PR_add[3][6] ), .OUT(m1614) );
  NOR2 U2538 ( .A(\PR_mul[5][7] ), .B(\PR_add[3][7] ), .OUT(m1615) );
  NOR2 U2539 ( .A(\PR_mul[5][8] ), .B(\PR_add[3][8] ), .OUT(m1616) );
  NOR2 U2540 ( .A(\PR_mul[5][9] ), .B(\PR_add[3][9] ), .OUT(m1617) );
  NOR2 U2541 ( .A(\PR_mul[5][10] ), .B(\PR_add[3][10] ), .OUT(m1618) );
  NAND2 U2542 ( .A(m1620), .B(\PR_add[3][18] ), .OUT(m1619) );
  NAND2 U2543 ( .A(\PR_add[3][15] ), .B(m1622), .OUT(m1621) );
  NOR2 U2544 ( .A(m1624), .B(m1625), .OUT(m1623) );
  NAND2 U2545 ( .A(m1627), .B(\PR_add[3][11] ), .OUT(m1626) );
  NOR2 U2546 ( .A(\PR_mul[4][3] ), .B(\PR_add[2][3] ), .OUT(m1628) );
  NOR2 U2547 ( .A(\PR_mul[4][4] ), .B(\PR_add[2][4] ), .OUT(m1629) );
  NOR2 U2548 ( .A(\PR_mul[4][5] ), .B(\PR_add[2][5] ), .OUT(m1630) );
  NOR2 U2549 ( .A(\PR_mul[4][6] ), .B(\PR_add[2][6] ), .OUT(m1631) );
  NOR2 U2550 ( .A(\PR_mul[4][7] ), .B(\PR_add[2][7] ), .OUT(m1632) );
  NOR2 U2551 ( .A(\PR_mul[4][8] ), .B(\PR_add[2][8] ), .OUT(m1633) );
  NOR2 U2552 ( .A(\PR_mul[4][9] ), .B(\PR_add[2][9] ), .OUT(m1634) );
  NOR2 U2553 ( .A(m1636), .B(m1637), .OUT(m1635) );
  NAND2 U2554 ( .A(\PR_add[2][16] ), .B(m1639), .OUT(m1638) );
  NAND2 U2555 ( .A(\PR_add[2][14] ), .B(m1641), .OUT(m1640) );
  NOR2 U2556 ( .A(m1643), .B(m1644), .OUT(m1642) );
  NAND2 U2557 ( .A(m1646), .B(\PR_add[2][10] ), .OUT(m1645) );
  NOR2 U2558 ( .A(\PR_mul[3][3] ), .B(\PR_add[1][3] ), .OUT(m1647) );
  NOR2 U2559 ( .A(\PR_mul[3][4] ), .B(\PR_add[1][4] ), .OUT(m1648) );
  NOR2 U2560 ( .A(\PR_mul[3][5] ), .B(\PR_add[1][5] ), .OUT(m1649) );
  NOR2 U2561 ( .A(\PR_mul[3][6] ), .B(\PR_add[1][6] ), .OUT(m1650) );
  NOR2 U2562 ( .A(\PR_mul[3][7] ), .B(\PR_add[1][7] ), .OUT(m1651) );
  NOR2 U2563 ( .A(\PR_mul[3][8] ), .B(\PR_add[1][8] ), .OUT(m1652) );
  NOR2 U2564 ( .A(\PR_mul[3][9] ), .B(\PR_add[1][9] ), .OUT(m1653) );
  NOR2 U2565 ( .A(\PR_mul[3][10] ), .B(\PR_add[1][10] ), .OUT(m1654) );
  NOR2 U2566 ( .A(\PR_mul[3][11] ), .B(\PR_add[1][11] ), .OUT(m1655) );
  NOR2 U2567 ( .A(m1657), .B(m1658), .OUT(m1656) );
  NAND2 U2568 ( .A(\PR_add[1][16] ), .B(m1660), .OUT(m1659) );
  NAND2 U2569 ( .A(m1662), .B(\PR_add[1][12] ), .OUT(m1661) );
  NOR2 U2570 ( .A(\PR_mul[2][1] ), .B(\PR_add[0][1] ), .OUT(m1663) );
  NOR2 U2571 ( .A(\PR_mul[2][2] ), .B(\PR_add[0][2] ), .OUT(m1664) );
  NOR2 U2572 ( .A(\PR_mul[2][3] ), .B(\PR_add[0][3] ), .OUT(m1665) );
  NOR2 U2573 ( .A(\PR_mul[2][4] ), .B(\PR_add[0][4] ), .OUT(m1666) );
  NOR2 U2574 ( .A(\PR_mul[2][5] ), .B(\PR_add[0][5] ), .OUT(m1667) );
  NOR2 U2575 ( .A(\PR_mul[2][6] ), .B(\PR_add[0][6] ), .OUT(m1668) );
  NOR2 U2576 ( .A(\PR_mul[2][7] ), .B(\PR_add[0][7] ), .OUT(m1669) );
  NOR2 U2577 ( .A(\PR_mul[2][8] ), .B(\PR_add[0][8] ), .OUT(m1670) );
  NOR2 U2578 ( .A(\PR_mul[2][9] ), .B(\PR_add[0][9] ), .OUT(m1671) );
  NOR2 U2579 ( .A(\PR_mul[2][10] ), .B(\PR_add[0][10] ), .OUT(m1672) );
  NOR2 U2580 ( .A(\PR_mul[2][11] ), .B(\PR_add[0][11] ), .OUT(m1673) );
  NOR2 U2581 ( .A(\PR_mul[1][4] ), .B(\PR_mul[0][4] ), .OUT(m1674) );
  NOR2 U2582 ( .A(\PR_mul[1][5] ), .B(\PR_mul[0][5] ), .OUT(m1675) );
  NOR2 U2583 ( .A(\PR_mul[1][6] ), .B(\PR_mul[0][6] ), .OUT(m1676) );
  NOR2 U2584 ( .A(\PR_mul[1][7] ), .B(\PR_mul[0][7] ), .OUT(m1677) );
  NOR2 U2585 ( .A(\PR_mul[1][8] ), .B(\PR_mul[0][8] ), .OUT(m1678) );
  NOR2 U2586 ( .A(\PR_mul[1][9] ), .B(\PR_mul[0][9] ), .OUT(m1679) );
  NOR2 U2587 ( .A(\PR_mul[1][10] ), .B(\PR_mul[0][10] ), .OUT(m1343) );
  XOR2 U2588 ( .A(m1339), .B(m1338), .OUT(\mult_83/A1[8] ) );
  XOR2 U2589 ( .A(m1680), .B(m1681), .OUT(\mult_83/A1[7] ) );
  XOR2 U2590 ( .A(m1682), .B(m1683), .OUT(\mult_83/A1[6] ) );
  XOR2 U2591 ( .A(m1684), .B(m1685), .OUT(\mult_83/A1[5] ) );
  XOR2 U2592 ( .A(m1686), .B(m1687), .OUT(\mult_83/A1[4] ) );
  XOR2 U2593 ( .A(m1688), .B(m1689), .OUT(\mult_83/A1[3] ) );
  XOR2 U2594 ( .A(m1317), .B(m1316), .OUT(\mult_82/A1[6] ) );
  XOR2 U2595 ( .A(m1690), .B(m1360), .OUT(\mult_82/A1[5] ) );
  XOR2 U2596 ( .A(m1691), .B(m1357), .OUT(\mult_82/A1[4] ) );
  XOR2 U2597 ( .A(m1692), .B(m1354), .OUT(\mult_82/A1[3] ) );
  XOR2 U2598 ( .A(\mult_80/ab[1][1] ), .B(\mult_80/ab[0][2] ), .OUT(m1693) );
  XOR2 U2599 ( .A(m1695), .B(m1696), .OUT(m1694) );
  XOR2 U2600 ( .A(m1335), .B(m1334), .OUT(\mult_80/A1[7] ) );
  XOR2 U2601 ( .A(m1694), .B(m1697), .OUT(\mult_80/A1[1] ) );
  XOR2 U2602 ( .A(m1333), .B(m1332), .OUT(\mult_77/A1[8] ) );
  XOR2 U2603 ( .A(m1698), .B(m1699), .OUT(\mult_77/A1[7] ) );
  XOR2 U2604 ( .A(m1700), .B(m1701), .OUT(\mult_77/A1[6] ) );
  XOR2 U2605 ( .A(m1702), .B(m1703), .OUT(\mult_77/A1[5] ) );
  XOR2 U2606 ( .A(m1704), .B(m1705), .OUT(\mult_77/A1[4] ) );
  XOR2 U2607 ( .A(m1706), .B(m1707), .OUT(\mult_77/A1[3] ) );
  XOR2 U2608 ( .A(m1331), .B(m1330), .OUT(\mult_76/A1[6] ) );
  XOR2 U2609 ( .A(m1708), .B(m1396), .OUT(\mult_76/A1[5] ) );
  XOR2 U2610 ( .A(m1709), .B(m1393), .OUT(\mult_76/A1[4] ) );
  XOR2 U2611 ( .A(m1710), .B(m1390), .OUT(\mult_76/A1[3] ) );
  XOR2 U2612 ( .A(\mult_74/ab[1][1] ), .B(\mult_74/ab[0][2] ), .OUT(m1711) );
  XOR2 U2613 ( .A(m1713), .B(m1714), .OUT(m1712) );
  XOR2 U2614 ( .A(m1327), .B(m1326), .OUT(\mult_74/A1[7] ) );
  XOR2 U2615 ( .A(m1712), .B(m1715), .OUT(\mult_74/A1[1] ) );
  XOR2 U2616 ( .A(m1325), .B(m1324), .OUT(\mult_72/A1[8] ) );
  XOR2 U2617 ( .A(m1716), .B(m1717), .OUT(\mult_72/A1[7] ) );
  XOR2 U2618 ( .A(m1718), .B(m1719), .OUT(\mult_72/A1[6] ) );
  XOR2 U2619 ( .A(m1720), .B(m1721), .OUT(\mult_72/A1[5] ) );
  XOR2 U2620 ( .A(m1722), .B(m1723), .OUT(\mult_72/A1[4] ) );
  XOR2 U2621 ( .A(m1724), .B(m1725), .OUT(\mult_72/A1[3] ) );
  XOR2 U2622 ( .A(m1323), .B(m1322), .OUT(\mult_71/A1[6] ) );
  XOR2 U2623 ( .A(m1726), .B(m1432), .OUT(\mult_71/A1[5] ) );
  XOR2 U2624 ( .A(m1727), .B(m1429), .OUT(\mult_71/A1[4] ) );
  XOR2 U2625 ( .A(m1728), .B(m1426), .OUT(\mult_71/A1[3] ) );
  XOR2 U2626 ( .A(\mult_69/ab[1][1] ), .B(\mult_69/ab[0][2] ), .OUT(m1729) );
  XOR2 U2627 ( .A(m1731), .B(m1732), .OUT(m1730) );
  XOR2 U2628 ( .A(m1319), .B(m1318), .OUT(\mult_69/A1[7] ) );
  XOR2 U2629 ( .A(m1730), .B(m1733), .OUT(\mult_69/A1[1] ) );
  XOR2 U2630 ( .A(\PR_add[12][10] ), .B(m1470), .OUT(N378) );
  XOR2 U2631 ( .A(m1734), .B(m1735), .OUT(N377) );
  XOR2 U2632 ( .A(m1736), .B(m1737), .OUT(N376) );
  XOR2 U2633 ( .A(m1738), .B(m1739), .OUT(N375) );
  XOR2 U2634 ( .A(m1740), .B(m1741), .OUT(N374) );
  XOR2 U2635 ( .A(m1742), .B(m1743), .OUT(N373) );
  XOR2 U2636 ( .A(m1744), .B(m1745), .OUT(N372) );
  XOR2 U2637 ( .A(\PR_add[11][12] ), .B(m1486), .OUT(N360) );
  XOR2 U2638 ( .A(m1746), .B(m1747), .OUT(N359) );
  XOR2 U2639 ( .A(m1748), .B(m1749), .OUT(N358) );
  XOR2 U2640 ( .A(m1750), .B(m1751), .OUT(N357) );
  XOR2 U2641 ( .A(m1752), .B(m1753), .OUT(N356) );
  XOR2 U2642 ( .A(m1754), .B(m1755), .OUT(N355) );
  XOR2 U2643 ( .A(m1756), .B(m1757), .OUT(N354) );
  XOR2 U2644 ( .A(m1758), .B(m1759), .OUT(N353) );
  XOR2 U2645 ( .A(m1760), .B(m1761), .OUT(N352) );
  XOR2 U2646 ( .A(m1762), .B(m1763), .OUT(N351) );
  XOR2 U2647 ( .A(\PR_add[10][12] ), .B(m1504), .OUT(N340) );
  XOR2 U2648 ( .A(m1764), .B(m1765), .OUT(N339) );
  XOR2 U2649 ( .A(m1766), .B(m1767), .OUT(N338) );
  XOR2 U2650 ( .A(m1768), .B(m1769), .OUT(N337) );
  XOR2 U2651 ( .A(m1770), .B(m1771), .OUT(N336) );
  XOR2 U2652 ( .A(m1772), .B(m1773), .OUT(N335) );
  XOR2 U2653 ( .A(m1774), .B(m1775), .OUT(N334) );
  XOR2 U2654 ( .A(m1776), .B(m1777), .OUT(N333) );
  XOR2 U2655 ( .A(m1778), .B(m1779), .OUT(N332) );
  XOR2 U2656 ( .A(m1780), .B(m1781), .OUT(N331) );
  XOR2 U2657 ( .A(m1782), .B(m1783), .OUT(N330) );
  XOR2 U2658 ( .A(\PR_add[9][11] ), .B(m1520), .OUT(N319) );
  XOR2 U2659 ( .A(m1784), .B(m1785), .OUT(N318) );
  XOR2 U2660 ( .A(m1786), .B(m1787), .OUT(N317) );
  XOR2 U2661 ( .A(m1788), .B(m1789), .OUT(N316) );
  XOR2 U2662 ( .A(m1790), .B(m1791), .OUT(N315) );
  XOR2 U2663 ( .A(m1792), .B(m1793), .OUT(N314) );
  XOR2 U2664 ( .A(m1794), .B(m1795), .OUT(N313) );
  XOR2 U2665 ( .A(\PR_add[8][11] ), .B(m1539), .OUT(N299) );
  XOR2 U2666 ( .A(m1796), .B(m1797), .OUT(N298) );
  XOR2 U2667 ( .A(m1798), .B(m1799), .OUT(N297) );
  XOR2 U2668 ( .A(m1800), .B(m1801), .OUT(N296) );
  XOR2 U2669 ( .A(m1802), .B(m1803), .OUT(N295) );
  XOR2 U2670 ( .A(m1804), .B(m1805), .OUT(N294) );
  XOR2 U2671 ( .A(m1806), .B(m1807), .OUT(N293) );
  XOR2 U2672 ( .A(m1808), .B(m1809), .OUT(N292) );
  XOR2 U2673 ( .A(m1810), .B(m1811), .OUT(N291) );
  XOR2 U2674 ( .A(m1812), .B(m1813), .OUT(N290) );
  XOR2 U2675 ( .A(\PR_add[7][10] ), .B(m1558), .OUT(N278) );
  XOR2 U2676 ( .A(m1814), .B(m1815), .OUT(N277) );
  XOR2 U2677 ( .A(m1816), .B(m1817), .OUT(N276) );
  XOR2 U2678 ( .A(m1818), .B(m1819), .OUT(N275) );
  XOR2 U2679 ( .A(m1820), .B(m1821), .OUT(N274) );
  XOR2 U2680 ( .A(m1822), .B(m1823), .OUT(N273) );
  XOR2 U2681 ( .A(m1824), .B(m1825), .OUT(N272) );
  XOR2 U2682 ( .A(\PR_add[6][12] ), .B(m1574), .OUT(N260) );
  XOR2 U2683 ( .A(m1826), .B(m1827), .OUT(N259) );
  XOR2 U2684 ( .A(m1828), .B(m1829), .OUT(N258) );
  XOR2 U2685 ( .A(m1830), .B(m1831), .OUT(N257) );
  XOR2 U2686 ( .A(m1832), .B(m1833), .OUT(N256) );
  XOR2 U2687 ( .A(m1834), .B(m1835), .OUT(N255) );
  XOR2 U2688 ( .A(m1836), .B(m1837), .OUT(N254) );
  XOR2 U2689 ( .A(m1838), .B(m1839), .OUT(N253) );
  XOR2 U2690 ( .A(m1840), .B(m1841), .OUT(N252) );
  XOR2 U2691 ( .A(m1842), .B(m1843), .OUT(N251) );
  XOR2 U2692 ( .A(\PR_add[5][12] ), .B(m1592), .OUT(N240) );
  XOR2 U2693 ( .A(m1844), .B(m1845), .OUT(N239) );
  XOR2 U2694 ( .A(m1846), .B(m1847), .OUT(N238) );
  XOR2 U2695 ( .A(m1848), .B(m1849), .OUT(N237) );
  XOR2 U2696 ( .A(m1850), .B(m1851), .OUT(N236) );
  XOR2 U2697 ( .A(m1852), .B(m1853), .OUT(N235) );
  XOR2 U2698 ( .A(m1854), .B(m1855), .OUT(N234) );
  XOR2 U2699 ( .A(m1856), .B(m1857), .OUT(N233) );
  XOR2 U2700 ( .A(m1858), .B(m1859), .OUT(N232) );
  XOR2 U2701 ( .A(m1860), .B(m1861), .OUT(N231) );
  XOR2 U2702 ( .A(m1862), .B(m1863), .OUT(N230) );
  XOR2 U2703 ( .A(\PR_add[4][11] ), .B(m1608), .OUT(N219) );
  XOR2 U2704 ( .A(m1864), .B(m1865), .OUT(N218) );
  XOR2 U2705 ( .A(m1866), .B(m1867), .OUT(N217) );
  XOR2 U2706 ( .A(m1868), .B(m1869), .OUT(N216) );
  XOR2 U2707 ( .A(m1870), .B(m1871), .OUT(N215) );
  XOR2 U2708 ( .A(m1872), .B(m1873), .OUT(N214) );
  XOR2 U2709 ( .A(m1874), .B(m1875), .OUT(N213) );
  XOR2 U2710 ( .A(\PR_add[3][11] ), .B(m1627), .OUT(N199) );
  XOR2 U2711 ( .A(m1876), .B(m1877), .OUT(N198) );
  XOR2 U2712 ( .A(m1878), .B(m1879), .OUT(N197) );
  XOR2 U2713 ( .A(m1880), .B(m1881), .OUT(N196) );
  XOR2 U2714 ( .A(m1882), .B(m1883), .OUT(N195) );
  XOR2 U2715 ( .A(m1884), .B(m1885), .OUT(N194) );
  XOR2 U2716 ( .A(m1886), .B(m1887), .OUT(N193) );
  XOR2 U2717 ( .A(m1888), .B(m1889), .OUT(N192) );
  XOR2 U2718 ( .A(m1890), .B(m1891), .OUT(N191) );
  XOR2 U2719 ( .A(m1892), .B(m1893), .OUT(N190) );
  XOR2 U2720 ( .A(\PR_add[2][10] ), .B(m1646), .OUT(N178) );
  XOR2 U2721 ( .A(m1894), .B(m1895), .OUT(N177) );
  XOR2 U2722 ( .A(m1896), .B(m1897), .OUT(N176) );
  XOR2 U2723 ( .A(m1898), .B(m1899), .OUT(N175) );
  XOR2 U2724 ( .A(m1900), .B(m1901), .OUT(N174) );
  XOR2 U2725 ( .A(m1902), .B(m1903), .OUT(N173) );
  XOR2 U2726 ( .A(m1904), .B(m1905), .OUT(N172) );
  XOR2 U2727 ( .A(\PR_add[1][12] ), .B(m1662), .OUT(N160) );
  XOR2 U2728 ( .A(m1906), .B(m1907), .OUT(N159) );
  XOR2 U2729 ( .A(m1908), .B(m1909), .OUT(N158) );
  XOR2 U2730 ( .A(m1910), .B(m1911), .OUT(N157) );
  XOR2 U2731 ( .A(m1912), .B(m1913), .OUT(N156) );
  XOR2 U2732 ( .A(m1914), .B(m1915), .OUT(N155) );
  XOR2 U2733 ( .A(m1916), .B(m1917), .OUT(N154) );
  XOR2 U2734 ( .A(m1918), .B(m1919), .OUT(N153) );
  XOR2 U2735 ( .A(m1920), .B(m1921), .OUT(N152) );
  XOR2 U2736 ( .A(m1922), .B(m1923), .OUT(N151) );
  XOR2 U2737 ( .A(m1924), .B(m1925), .OUT(N139) );
  XOR2 U2738 ( .A(m1926), .B(m1927), .OUT(N138) );
  XOR2 U2739 ( .A(m1928), .B(m1929), .OUT(N137) );
  XOR2 U2740 ( .A(m1930), .B(m1931), .OUT(N136) );
  XOR2 U2741 ( .A(m1932), .B(m1933), .OUT(N135) );
  XOR2 U2742 ( .A(m1934), .B(m1935), .OUT(N134) );
  XOR2 U2743 ( .A(m1936), .B(m1937), .OUT(N133) );
  XOR2 U2744 ( .A(m1938), .B(m1939), .OUT(N132) );
  XOR2 U2745 ( .A(m1940), .B(m1941), .OUT(N131) );
  XOR2 U2746 ( .A(m1942), .B(m1943), .OUT(N130) );
  XOR2 U2747 ( .A(m1944), .B(m1342), .OUT(N118) );
  XOR2 U2748 ( .A(m1945), .B(m1946), .OUT(N117) );
  XOR2 U2749 ( .A(m1947), .B(m1948), .OUT(N116) );
  XOR2 U2750 ( .A(m1949), .B(m1950), .OUT(N115) );
  XOR2 U2751 ( .A(m1951), .B(m1952), .OUT(N114) );
  XOR2 U2752 ( .A(m1953), .B(m1954), .OUT(N113) );
  NAND2 U2753 ( .A(\mult_83/ab[0][3] ), .B(\mult_83/ab[1][2] ), .OUT(m1955) );
  INV U2754 ( .IN(\mult_83/ab[7][3] ), .OUT(m1339) );
  NAND2 U2755 ( .A(\mult_82/ab[0][3] ), .B(\mult_82/ab[3][0] ), .OUT(m1956) );
  AOI22 U2756 ( .A(\mult_82/ab[4][0] ), .B(m1351), .C(m1957), .D(
        \mult_82/ab[1][3] ), .OUT(m1354) );
  INV U2757 ( .IN(\mult_82/ab[5][0] ), .OUT(m1353) );
  AOI22 U2758 ( .A(m1958), .B(\mult_82/ab[5][0] ), .C(m1352), .D(
        \mult_82/ab[2][3] ), .OUT(m1357) );
  INV U2759 ( .IN(\mult_82/ab[6][0] ), .OUT(m1356) );
  AOI22 U2760 ( .A(m1959), .B(\mult_82/ab[6][0] ), .C(m1355), .D(
        \mult_82/ab[3][3] ), .OUT(m1360) );
  INV U2761 ( .IN(\mult_82/ab[7][0] ), .OUT(m1359) );
  INV U2762 ( .IN(\mult_82/ab[5][3] ), .OUT(m1317) );
  NAND2 U2763 ( .A(\mult_80/ab[0][2] ), .B(\mult_80/ab[1][1] ), .OUT(m1960) );
  INV U2764 ( .IN(\mult_80/ab[1][2] ), .OUT(m1695) );
  INV U2765 ( .IN(\mult_80/ab[2][1] ), .OUT(m1961) );
  INV U2766 ( .IN(\mult_80/ab[7][2] ), .OUT(m1335) );
  NAND2 U2767 ( .A(\mult_80/ab[0][1] ), .B(\mult_80/ab[1][0] ), .OUT(m1369) );
  AOI22 U2768 ( .A(\mult_80/ab[2][0] ), .B(m1963), .C(m1367), .D(m1693), .OUT(
        m1962) );
  INV U2769 ( .IN(\mult_80/ab[3][0] ), .OUT(m1964) );
  OAI22 U2770 ( .A(m1962), .B(m1964), .C(m1370), .D(m1694), .OUT(m1373) );
  AOI22 U2771 ( .A(m1373), .B(\mult_80/ab[4][0] ), .C(m1966), .D(m1967), .OUT(
        m1965) );
  INV U2772 ( .IN(\mult_80/ab[5][0] ), .OUT(m1968) );
  OAI22 U2773 ( .A(m1965), .B(m1968), .C(m1374), .D(m1969), .OUT(m1377) );
  INV U2774 ( .IN(\mult_80/ab[6][0] ), .OUT(m1970) );
  OAI22 U2775 ( .A(m1971), .B(m1970), .C(m1376), .D(m1972), .OUT(m1379) );
  NAND2 U2776 ( .A(\mult_77/ab[0][3] ), .B(\mult_77/ab[1][2] ), .OUT(m1973) );
  INV U2777 ( .IN(\mult_77/ab[7][3] ), .OUT(m1333) );
  NAND2 U2778 ( .A(\mult_76/ab[0][3] ), .B(\mult_76/ab[3][0] ), .OUT(m1974) );
  AOI22 U2779 ( .A(\mult_76/ab[4][0] ), .B(m1387), .C(m1975), .D(
        \mult_76/ab[1][3] ), .OUT(m1390) );
  INV U2780 ( .IN(\mult_76/ab[5][0] ), .OUT(m1389) );
  AOI22 U2781 ( .A(m1976), .B(\mult_76/ab[5][0] ), .C(m1388), .D(
        \mult_76/ab[2][3] ), .OUT(m1393) );
  INV U2782 ( .IN(\mult_76/ab[6][0] ), .OUT(m1392) );
  AOI22 U2783 ( .A(m1977), .B(\mult_76/ab[6][0] ), .C(m1391), .D(
        \mult_76/ab[3][3] ), .OUT(m1396) );
  INV U2784 ( .IN(\mult_76/ab[7][0] ), .OUT(m1395) );
  INV U2785 ( .IN(\mult_76/ab[5][3] ), .OUT(m1331) );
  NAND2 U2786 ( .A(\mult_74/ab[0][2] ), .B(\mult_74/ab[1][1] ), .OUT(m1978) );
  INV U2787 ( .IN(\mult_74/ab[1][2] ), .OUT(m1713) );
  INV U2788 ( .IN(\mult_74/ab[2][1] ), .OUT(m1979) );
  INV U2789 ( .IN(\mult_74/ab[7][2] ), .OUT(m1327) );
  NAND2 U2790 ( .A(\mult_74/ab[0][1] ), .B(\mult_74/ab[1][0] ), .OUT(m1405) );
  AOI22 U2791 ( .A(\mult_74/ab[2][0] ), .B(m1981), .C(m1403), .D(m1711), .OUT(
        m1980) );
  INV U2792 ( .IN(\mult_74/ab[3][0] ), .OUT(m1982) );
  OAI22 U2793 ( .A(m1980), .B(m1982), .C(m1406), .D(m1712), .OUT(m1409) );
  AOI22 U2794 ( .A(m1409), .B(\mult_74/ab[4][0] ), .C(m1984), .D(m1985), .OUT(
        m1983) );
  INV U2795 ( .IN(\mult_74/ab[5][0] ), .OUT(m1986) );
  OAI22 U2796 ( .A(m1983), .B(m1986), .C(m1410), .D(m1987), .OUT(m1413) );
  INV U2797 ( .IN(\mult_74/ab[6][0] ), .OUT(m1988) );
  OAI22 U2798 ( .A(m1989), .B(m1988), .C(m1412), .D(m1990), .OUT(m1415) );
  NAND2 U2799 ( .A(\mult_72/ab[0][3] ), .B(\mult_72/ab[1][2] ), .OUT(m1991) );
  INV U2800 ( .IN(\mult_72/ab[7][3] ), .OUT(m1325) );
  NAND2 U2801 ( .A(\mult_71/ab[0][3] ), .B(\mult_71/ab[3][0] ), .OUT(m1992) );
  AOI22 U2802 ( .A(\mult_71/ab[4][0] ), .B(m1423), .C(m1993), .D(
        \mult_71/ab[1][3] ), .OUT(m1426) );
  INV U2803 ( .IN(\mult_71/ab[5][0] ), .OUT(m1425) );
  AOI22 U2804 ( .A(m1994), .B(\mult_71/ab[5][0] ), .C(m1424), .D(
        \mult_71/ab[2][3] ), .OUT(m1429) );
  INV U2805 ( .IN(\mult_71/ab[6][0] ), .OUT(m1428) );
  AOI22 U2806 ( .A(m1995), .B(\mult_71/ab[6][0] ), .C(m1427), .D(
        \mult_71/ab[3][3] ), .OUT(m1432) );
  INV U2807 ( .IN(\mult_71/ab[7][0] ), .OUT(m1431) );
  INV U2808 ( .IN(\mult_71/ab[5][3] ), .OUT(m1323) );
  NAND2 U2809 ( .A(\mult_69/ab[0][2] ), .B(\mult_69/ab[1][1] ), .OUT(m1996) );
  INV U2810 ( .IN(\mult_69/ab[1][2] ), .OUT(m1731) );
  INV U2811 ( .IN(\mult_69/ab[2][1] ), .OUT(m1997) );
  INV U2812 ( .IN(\mult_69/ab[7][2] ), .OUT(m1319) );
  NAND2 U2813 ( .A(\mult_69/ab[0][1] ), .B(\mult_69/ab[1][0] ), .OUT(m1441) );
  AOI22 U2814 ( .A(\mult_69/ab[2][0] ), .B(m1999), .C(m1439), .D(m1729), .OUT(
        m1998) );
  INV U2815 ( .IN(\mult_69/ab[3][0] ), .OUT(m2000) );
  OAI22 U2816 ( .A(m1998), .B(m2000), .C(m1442), .D(m1730), .OUT(m1445) );
  AOI22 U2817 ( .A(m1445), .B(\mult_69/ab[4][0] ), .C(m2002), .D(m2003), .OUT(
        m2001) );
  INV U2818 ( .IN(\mult_69/ab[5][0] ), .OUT(m2004) );
  OAI22 U2819 ( .A(m2001), .B(m2004), .C(m1446), .D(m2005), .OUT(m1449) );
  INV U2820 ( .IN(\mult_69/ab[6][0] ), .OUT(m2006) );
  OAI22 U2821 ( .A(m2007), .B(m2006), .C(m1448), .D(m2008), .OUT(m1451) );
  NAND2 U2822 ( .A(\PR_add[12][2] ), .B(\PR_mul[14][2] ), .OUT(m2009) );
  INV U2823 ( .IN(\PR_mul[14][9] ), .OUT(m2010) );
  INV U2824 ( .IN(\PR_add[12][9] ), .OUT(m2011) );
  INV U2825 ( .IN(\PR_add[12][12] ), .OUT(m1467) );
  NAND3 U2826 ( .A(\PR_add[12][11] ), .B(m1470), .C(\PR_add[12][10] ), .OUT(
        m1468) );
  NOR3 U2827 ( .A(m1467), .B(m2012), .C(m1468), .OUT(m1465) );
  NAND3 U2828 ( .A(\PR_add[12][14] ), .B(\PR_add[12][15] ), .C(m1465), .OUT(
        m2013) );
  INV U2829 ( .IN(\PR_add[12][18] ), .OUT(m1460) );
  NAND3 U2830 ( .A(\PR_add[12][16] ), .B(\PR_add[12][17] ), .C(m1463), .OUT(
        m1461) );
  INV U2831 ( .IN(\PR_mul[13][11] ), .OUT(m2015) );
  INV U2832 ( .IN(\PR_add[11][11] ), .OUT(m2016) );
  INV U2833 ( .IN(\PR_add[11][15] ), .OUT(m2017) );
  INV U2834 ( .IN(\PR_add[11][14] ), .OUT(m2018) );
  NAND3 U2835 ( .A(\PR_add[11][13] ), .B(m1486), .C(\PR_add[11][12] ), .OUT(
        m2019) );
  NOR3 U2836 ( .A(m2018), .B(m2017), .C(m2019), .OUT(m1484) );
  INV U2837 ( .IN(\PR_add[11][18] ), .OUT(m1481) );
  NAND3 U2838 ( .A(\PR_add[11][16] ), .B(\PR_add[11][17] ), .C(m1484), .OUT(
        m1482) );
  NAND2 U2839 ( .A(\PR_add[10][0] ), .B(\PR_mul[12][0] ), .OUT(m2020) );
  INV U2840 ( .IN(\PR_mul[12][11] ), .OUT(m2021) );
  INV U2841 ( .IN(\PR_add[10][11] ), .OUT(m2022) );
  INV U2842 ( .IN(\PR_add[10][15] ), .OUT(m2023) );
  INV U2843 ( .IN(\PR_add[10][14] ), .OUT(m2024) );
  NAND3 U2844 ( .A(\PR_add[10][13] ), .B(m1504), .C(\PR_add[10][12] ), .OUT(
        m2025) );
  NOR3 U2845 ( .A(m2024), .B(m2023), .C(m2025), .OUT(m1502) );
  INV U2846 ( .IN(\PR_add[10][18] ), .OUT(m1499) );
  NAND3 U2847 ( .A(\PR_add[10][16] ), .B(\PR_add[10][17] ), .C(m1502), .OUT(
        m1500) );
  NAND2 U2848 ( .A(\PR_add[9][3] ), .B(\PR_mul[11][3] ), .OUT(m2026) );
  INV U2849 ( .IN(\PR_mul[11][10] ), .OUT(m2027) );
  INV U2850 ( .IN(\PR_add[9][10] ), .OUT(m2028) );
  INV U2851 ( .IN(\PR_add[9][13] ), .OUT(m1517) );
  NAND3 U2852 ( .A(\PR_add[9][12] ), .B(m1520), .C(\PR_add[9][11] ), .OUT(
        m1518) );
  NOR3 U2853 ( .A(m1517), .B(m2029), .C(m1518), .OUT(m1515) );
  INV U2854 ( .IN(\PR_add[9][17] ), .OUT(m2030) );
  NAND3 U2855 ( .A(\PR_add[9][15] ), .B(\PR_add[9][16] ), .C(m1515), .OUT(
        m2031) );
  NOR2 U2856 ( .A(m2031), .B(m2030), .OUT(m1513) );
  NAND2 U2857 ( .A(\PR_add[8][0] ), .B(\PR_mul[10][0] ), .OUT(m2032) );
  INV U2858 ( .IN(\PR_mul[10][10] ), .OUT(m2033) );
  INV U2859 ( .IN(\PR_add[8][10] ), .OUT(m2034) );
  INV U2860 ( .IN(\PR_add[8][13] ), .OUT(m1536) );
  NAND3 U2861 ( .A(\PR_add[8][12] ), .B(m1539), .C(\PR_add[8][11] ), .OUT(
        m1537) );
  NOR3 U2862 ( .A(m1536), .B(m2035), .C(m1537), .OUT(m1534) );
  INV U2863 ( .IN(\PR_add[8][17] ), .OUT(m2036) );
  NAND3 U2864 ( .A(\PR_add[8][15] ), .B(\PR_add[8][16] ), .C(m1534), .OUT(
        m2037) );
  NOR2 U2865 ( .A(m2037), .B(m2036), .OUT(m1532) );
  NAND2 U2866 ( .A(\PR_add[7][2] ), .B(\PR_mul[9][2] ), .OUT(m2038) );
  INV U2867 ( .IN(\PR_mul[9][9] ), .OUT(m2039) );
  INV U2868 ( .IN(\PR_add[7][9] ), .OUT(m2040) );
  INV U2869 ( .IN(\PR_add[7][12] ), .OUT(m1555) );
  NAND3 U2870 ( .A(\PR_add[7][11] ), .B(m1558), .C(\PR_add[7][10] ), .OUT(
        m1556) );
  NOR3 U2871 ( .A(m1555), .B(m2041), .C(m1556), .OUT(m1553) );
  NAND3 U2872 ( .A(\PR_add[7][14] ), .B(\PR_add[7][15] ), .C(m1553), .OUT(
        m2042) );
  INV U2873 ( .IN(\PR_add[7][18] ), .OUT(m1548) );
  NAND3 U2874 ( .A(\PR_add[7][16] ), .B(\PR_add[7][17] ), .C(m1551), .OUT(
        m1549) );
  INV U2875 ( .IN(\PR_mul[8][11] ), .OUT(m2044) );
  INV U2876 ( .IN(\PR_add[6][11] ), .OUT(m2045) );
  INV U2877 ( .IN(\PR_add[6][15] ), .OUT(m2046) );
  INV U2878 ( .IN(\PR_add[6][14] ), .OUT(m2047) );
  NAND3 U2879 ( .A(\PR_add[6][13] ), .B(m1574), .C(\PR_add[6][12] ), .OUT(
        m2048) );
  NOR3 U2880 ( .A(m2047), .B(m2046), .C(m2048), .OUT(m1572) );
  INV U2881 ( .IN(\PR_add[6][18] ), .OUT(m1569) );
  NAND3 U2882 ( .A(\PR_add[6][16] ), .B(\PR_add[6][17] ), .C(m1572), .OUT(
        m1570) );
  NAND2 U2883 ( .A(\PR_add[5][0] ), .B(\PR_mul[7][0] ), .OUT(m2049) );
  INV U2884 ( .IN(\PR_mul[7][11] ), .OUT(m2050) );
  INV U2885 ( .IN(\PR_add[5][11] ), .OUT(m2051) );
  INV U2886 ( .IN(\PR_add[5][15] ), .OUT(m2052) );
  INV U2887 ( .IN(\PR_add[5][14] ), .OUT(m2053) );
  NAND3 U2888 ( .A(\PR_add[5][13] ), .B(m1592), .C(\PR_add[5][12] ), .OUT(
        m2054) );
  NOR3 U2889 ( .A(m2053), .B(m2052), .C(m2054), .OUT(m1590) );
  INV U2890 ( .IN(\PR_add[5][18] ), .OUT(m1587) );
  NAND3 U2891 ( .A(\PR_add[5][16] ), .B(\PR_add[5][17] ), .C(m1590), .OUT(
        m1588) );
  NAND2 U2892 ( .A(\PR_add[4][3] ), .B(\PR_mul[6][3] ), .OUT(m2055) );
  INV U2893 ( .IN(\PR_mul[6][10] ), .OUT(m2056) );
  INV U2894 ( .IN(\PR_add[4][10] ), .OUT(m2057) );
  INV U2895 ( .IN(\PR_add[4][13] ), .OUT(m1605) );
  NAND3 U2896 ( .A(\PR_add[4][12] ), .B(m1608), .C(\PR_add[4][11] ), .OUT(
        m1606) );
  NOR3 U2897 ( .A(m1605), .B(m2058), .C(m1606), .OUT(m1603) );
  INV U2898 ( .IN(\PR_add[4][17] ), .OUT(m2059) );
  NAND3 U2899 ( .A(\PR_add[4][15] ), .B(\PR_add[4][16] ), .C(m1603), .OUT(
        m2060) );
  NOR2 U2900 ( .A(m2060), .B(m2059), .OUT(m1601) );
  NAND2 U2901 ( .A(\PR_add[3][0] ), .B(\PR_mul[5][0] ), .OUT(m2061) );
  INV U2902 ( .IN(\PR_mul[5][10] ), .OUT(m2062) );
  INV U2903 ( .IN(\PR_add[3][10] ), .OUT(m2063) );
  INV U2904 ( .IN(\PR_add[3][13] ), .OUT(m1624) );
  NAND3 U2905 ( .A(\PR_add[3][12] ), .B(m1627), .C(\PR_add[3][11] ), .OUT(
        m1625) );
  NOR3 U2906 ( .A(m1624), .B(m2064), .C(m1625), .OUT(m1622) );
  INV U2907 ( .IN(\PR_add[3][17] ), .OUT(m2065) );
  NAND3 U2908 ( .A(\PR_add[3][15] ), .B(\PR_add[3][16] ), .C(m1622), .OUT(
        m2066) );
  NOR2 U2909 ( .A(m2066), .B(m2065), .OUT(m1620) );
  NAND2 U2910 ( .A(\PR_add[2][2] ), .B(\PR_mul[4][2] ), .OUT(m2067) );
  INV U2911 ( .IN(\PR_mul[4][9] ), .OUT(m2068) );
  INV U2912 ( .IN(\PR_add[2][9] ), .OUT(m2069) );
  INV U2913 ( .IN(\PR_add[2][12] ), .OUT(m1643) );
  NAND3 U2914 ( .A(\PR_add[2][11] ), .B(m1646), .C(\PR_add[2][10] ), .OUT(
        m1644) );
  NOR3 U2915 ( .A(m1643), .B(m2070), .C(m1644), .OUT(m1641) );
  NAND3 U2916 ( .A(\PR_add[2][14] ), .B(\PR_add[2][15] ), .C(m1641), .OUT(
        m2071) );
  INV U2917 ( .IN(\PR_add[2][18] ), .OUT(m1636) );
  NAND3 U2918 ( .A(\PR_add[2][16] ), .B(\PR_add[2][17] ), .C(m1639), .OUT(
        m1637) );
  INV U2919 ( .IN(\PR_mul[3][11] ), .OUT(m2073) );
  INV U2920 ( .IN(\PR_add[1][11] ), .OUT(m2074) );
  INV U2921 ( .IN(\PR_add[1][15] ), .OUT(m2075) );
  INV U2922 ( .IN(\PR_add[1][14] ), .OUT(m2076) );
  NAND3 U2923 ( .A(\PR_add[1][13] ), .B(m1662), .C(\PR_add[1][12] ), .OUT(
        m2077) );
  NOR3 U2924 ( .A(m2076), .B(m2075), .C(m2077), .OUT(m1660) );
  INV U2925 ( .IN(\PR_add[1][18] ), .OUT(m1657) );
  NAND3 U2926 ( .A(\PR_add[1][16] ), .B(\PR_add[1][17] ), .C(m1660), .OUT(
        m1658) );
  NAND2 U2927 ( .A(\PR_add[0][0] ), .B(\PR_mul[2][0] ), .OUT(m2078) );
  INV U2928 ( .IN(\PR_mul[2][11] ), .OUT(m2079) );
  INV U2929 ( .IN(\PR_add[0][11] ), .OUT(m2080) );
  NAND2 U2930 ( .A(\PR_mul[0][3] ), .B(\PR_mul[1][3] ), .OUT(m2081) );
  INV U2931 ( .IN(\PR_mul[1][10] ), .OUT(m1340) );
  INV U2932 ( .IN(\PR_mul[0][10] ), .OUT(m1341) );
  XOR2 U2933 ( .A(m2082), .B(m2083), .OUT(\mult_83/A1[2] ) );
  XOR2 U2934 ( .A(\mult_83/ab[0][3] ), .B(\mult_83/ab[1][2] ), .OUT(
        \mult_83/A1[1] ) );
  XOR2 U2935 ( .A(\mult_82/ab[4][0] ), .B(m2084), .OUT(\mult_82/A1[2] ) );
  XOR2 U2936 ( .A(\mult_82/ab[0][3] ), .B(\mult_82/ab[3][0] ), .OUT(
        \mult_82/A1[1] ) );
  XOR2 U2937 ( .A(m1336), .B(m1337), .OUT(\mult_80/A1[6] ) );
  XOR2 U2938 ( .A(m2085), .B(m2086), .OUT(\mult_80/A1[5] ) );
  XOR2 U2939 ( .A(m1972), .B(m2087), .OUT(\mult_80/A1[4] ) );
  XOR2 U2940 ( .A(m1969), .B(m2088), .OUT(\mult_80/A1[3] ) );
  XOR2 U2941 ( .A(m1967), .B(m2089), .OUT(\mult_80/A1[2] ) );
  XOR2 U2942 ( .A(m1693), .B(m2090), .OUT(\mult_80/A1[0] ) );
  XOR2 U2943 ( .A(m2091), .B(m2092), .OUT(\mult_77/A1[2] ) );
  XOR2 U2944 ( .A(\mult_77/ab[0][3] ), .B(\mult_77/ab[1][2] ), .OUT(
        \mult_77/A1[1] ) );
  XOR2 U2945 ( .A(\mult_76/ab[4][0] ), .B(m2093), .OUT(\mult_76/A1[2] ) );
  XOR2 U2946 ( .A(\mult_76/ab[0][3] ), .B(\mult_76/ab[3][0] ), .OUT(
        \mult_76/A1[1] ) );
  XOR2 U2947 ( .A(m1328), .B(m1329), .OUT(\mult_74/A1[6] ) );
  XOR2 U2948 ( .A(m2094), .B(m2095), .OUT(\mult_74/A1[5] ) );
  XOR2 U2949 ( .A(m1990), .B(m2096), .OUT(\mult_74/A1[4] ) );
  XOR2 U2950 ( .A(m1987), .B(m2097), .OUT(\mult_74/A1[3] ) );
  XOR2 U2951 ( .A(m1985), .B(m2098), .OUT(\mult_74/A1[2] ) );
  XOR2 U2952 ( .A(m1711), .B(m2099), .OUT(\mult_74/A1[0] ) );
  XOR2 U2953 ( .A(m2100), .B(m2101), .OUT(\mult_72/A1[2] ) );
  XOR2 U2954 ( .A(\mult_72/ab[0][3] ), .B(\mult_72/ab[1][2] ), .OUT(
        \mult_72/A1[1] ) );
  XOR2 U2955 ( .A(\mult_71/ab[4][0] ), .B(m2102), .OUT(\mult_71/A1[2] ) );
  XOR2 U2956 ( .A(\mult_71/ab[0][3] ), .B(\mult_71/ab[3][0] ), .OUT(
        \mult_71/A1[1] ) );
  XOR2 U2957 ( .A(m1320), .B(m1321), .OUT(\mult_69/A1[6] ) );
  XOR2 U2958 ( .A(m2103), .B(m2104), .OUT(\mult_69/A1[5] ) );
  XOR2 U2959 ( .A(m2008), .B(m2105), .OUT(\mult_69/A1[4] ) );
  XOR2 U2960 ( .A(m2005), .B(m2106), .OUT(\mult_69/A1[3] ) );
  XOR2 U2961 ( .A(m2003), .B(m2107), .OUT(\mult_69/A1[2] ) );
  XOR2 U2962 ( .A(m1729), .B(m2108), .OUT(\mult_69/A1[0] ) );
  XOR2 U2963 ( .A(\mult_80/ab[0][1] ), .B(\mult_80/ab[1][0] ), .OUT(N74) );
  XOR2 U2964 ( .A(\mult_69/ab[0][1] ), .B(\mult_69/ab[1][0] ), .OUT(N4) );
  XOR2 U2965 ( .A(\mult_74/ab[0][1] ), .B(\mult_74/ab[1][0] ), .OUT(N39) );
  XOR2 U2966 ( .A(\PR_add[12][19] ), .B(m1459), .OUT(N387) );
  XOR2 U2967 ( .A(m1461), .B(m1460), .OUT(N386) );
  XOR2 U2968 ( .A(\PR_add[12][17] ), .B(m1462), .OUT(m2109) );
  XOR2 U2969 ( .A(m1463), .B(\PR_add[12][16] ), .OUT(N384) );
  XOR2 U2970 ( .A(\PR_add[12][15] ), .B(m1464), .OUT(m2110) );
  XOR2 U2971 ( .A(m1465), .B(\PR_add[12][14] ), .OUT(N382) );
  XOR2 U2972 ( .A(\PR_add[12][13] ), .B(m1466), .OUT(N381) );
  XOR2 U2973 ( .A(m1468), .B(m1467), .OUT(N380) );
  XOR2 U2974 ( .A(\PR_add[12][11] ), .B(m1469), .OUT(m2111) );
  XOR2 U2975 ( .A(m2112), .B(m2113), .OUT(N371) );
  XOR2 U2976 ( .A(\PR_add[12][2] ), .B(\PR_mul[14][2] ), .OUT(N370) );
  XOR2 U2977 ( .A(\PR_add[11][19] ), .B(m1480), .OUT(N367) );
  XOR2 U2978 ( .A(m1482), .B(m1481), .OUT(N366) );
  XOR2 U2979 ( .A(\PR_add[11][17] ), .B(m1483), .OUT(m2114) );
  XOR2 U2980 ( .A(m1484), .B(\PR_add[11][16] ), .OUT(N364) );
  XOR2 U2981 ( .A(\PR_add[11][15] ), .B(m2115), .OUT(N363) );
  XOR2 U2982 ( .A(m2019), .B(m2018), .OUT(N362) );
  XOR2 U2983 ( .A(\PR_add[11][13] ), .B(m1485), .OUT(m2116) );
  XOR2 U2984 ( .A(\PR_add[10][19] ), .B(m1498), .OUT(N347) );
  XOR2 U2985 ( .A(m1500), .B(m1499), .OUT(N346) );
  XOR2 U2986 ( .A(\PR_add[10][17] ), .B(m1501), .OUT(m2119) );
  XOR2 U2987 ( .A(m1502), .B(\PR_add[10][16] ), .OUT(N344) );
  XOR2 U2988 ( .A(\PR_add[10][15] ), .B(m2120), .OUT(N343) );
  XOR2 U2989 ( .A(m2025), .B(m2024), .OUT(N342) );
  XOR2 U2990 ( .A(\PR_add[10][13] ), .B(m1503), .OUT(m2121) );
  XOR2 U2991 ( .A(m2122), .B(m2123), .OUT(N329) );
  XOR2 U2992 ( .A(\PR_add[10][0] ), .B(\PR_mul[12][0] ), .OUT(N328) );
  XOR2 U2993 ( .A(\PR_add[9][19] ), .B(m1512), .OUT(m2124) );
  XOR2 U2994 ( .A(\PR_add[9][18] ), .B(m1513), .OUT(N326) );
  XOR2 U2995 ( .A(m2031), .B(m2030), .OUT(N325) );
  XOR2 U2996 ( .A(\PR_add[9][16] ), .B(m1514), .OUT(m2125) );
  XOR2 U2997 ( .A(m1515), .B(\PR_add[9][15] ), .OUT(N323) );
  XOR2 U2998 ( .A(\PR_add[9][14] ), .B(m1516), .OUT(N322) );
  XOR2 U2999 ( .A(m1518), .B(m1517), .OUT(N321) );
  XOR2 U3000 ( .A(\PR_add[9][12] ), .B(m1519), .OUT(m2126) );
  XOR2 U3001 ( .A(m2127), .B(m2128), .OUT(N312) );
  XOR2 U3002 ( .A(\PR_add[9][3] ), .B(\PR_mul[11][3] ), .OUT(N311) );
  XOR2 U3003 ( .A(\PR_add[8][19] ), .B(m1531), .OUT(m2129) );
  XOR2 U3004 ( .A(\PR_add[8][18] ), .B(m1532), .OUT(N306) );
  XOR2 U3005 ( .A(m2037), .B(m2036), .OUT(N305) );
  XOR2 U3006 ( .A(\PR_add[8][16] ), .B(m1533), .OUT(m2130) );
  XOR2 U3007 ( .A(m1534), .B(\PR_add[8][15] ), .OUT(N303) );
  XOR2 U3008 ( .A(\PR_add[8][14] ), .B(m1535), .OUT(N302) );
  XOR2 U3009 ( .A(m1537), .B(m1536), .OUT(N301) );
  XOR2 U3010 ( .A(\PR_add[8][12] ), .B(m1538), .OUT(m2131) );
  XOR2 U3011 ( .A(m2132), .B(m2133), .OUT(N289) );
  XOR2 U3012 ( .A(\PR_add[8][0] ), .B(\PR_mul[10][0] ), .OUT(N288) );
  XOR2 U3013 ( .A(\PR_add[7][19] ), .B(m1547), .OUT(N287) );
  XOR2 U3014 ( .A(m1549), .B(m1548), .OUT(N286) );
  XOR2 U3015 ( .A(\PR_add[7][17] ), .B(m1550), .OUT(m2134) );
  XOR2 U3016 ( .A(m1551), .B(\PR_add[7][16] ), .OUT(N284) );
  XOR2 U3017 ( .A(\PR_add[7][15] ), .B(m1552), .OUT(m2135) );
  XOR2 U3018 ( .A(m1553), .B(\PR_add[7][14] ), .OUT(N282) );
  XOR2 U3019 ( .A(\PR_add[7][13] ), .B(m1554), .OUT(N281) );
  XOR2 U3020 ( .A(m1556), .B(m1555), .OUT(N280) );
  XOR2 U3021 ( .A(\PR_add[7][11] ), .B(m1557), .OUT(m2136) );
  XOR2 U3022 ( .A(m2137), .B(m2138), .OUT(N271) );
  XOR2 U3023 ( .A(\PR_add[7][2] ), .B(\PR_mul[9][2] ), .OUT(N270) );
  XOR2 U3024 ( .A(\PR_add[6][19] ), .B(m1568), .OUT(N267) );
  XOR2 U3025 ( .A(m1570), .B(m1569), .OUT(N266) );
  XOR2 U3026 ( .A(\PR_add[6][17] ), .B(m1571), .OUT(m2139) );
  XOR2 U3027 ( .A(m1572), .B(\PR_add[6][16] ), .OUT(N264) );
  XOR2 U3028 ( .A(\PR_add[6][15] ), .B(m2140), .OUT(N263) );
  XOR2 U3029 ( .A(m2048), .B(m2047), .OUT(N262) );
  XOR2 U3030 ( .A(\PR_add[6][13] ), .B(m1573), .OUT(m2141) );
  XOR2 U3031 ( .A(\PR_add[5][19] ), .B(m1586), .OUT(N247) );
  XOR2 U3032 ( .A(m1588), .B(m1587), .OUT(N246) );
  XOR2 U3033 ( .A(\PR_add[5][17] ), .B(m1589), .OUT(m2144) );
  XOR2 U3034 ( .A(m1590), .B(\PR_add[5][16] ), .OUT(N244) );
  XOR2 U3035 ( .A(\PR_add[5][15] ), .B(m2145), .OUT(N243) );
  XOR2 U3036 ( .A(m2054), .B(m2053), .OUT(N242) );
  XOR2 U3037 ( .A(\PR_add[5][13] ), .B(m1591), .OUT(m2146) );
  XOR2 U3038 ( .A(m2147), .B(m2148), .OUT(N229) );
  XOR2 U3039 ( .A(\PR_add[5][0] ), .B(\PR_mul[7][0] ), .OUT(N228) );
  XOR2 U3040 ( .A(\PR_add[4][19] ), .B(m1600), .OUT(m2149) );
  XOR2 U3041 ( .A(\PR_add[4][18] ), .B(m1601), .OUT(N226) );
  XOR2 U3042 ( .A(m2060), .B(m2059), .OUT(N225) );
  XOR2 U3043 ( .A(\PR_add[4][16] ), .B(m1602), .OUT(m2150) );
  XOR2 U3044 ( .A(m1603), .B(\PR_add[4][15] ), .OUT(N223) );
  XOR2 U3045 ( .A(\PR_add[4][14] ), .B(m1604), .OUT(N222) );
  XOR2 U3046 ( .A(m1606), .B(m1605), .OUT(N221) );
  XOR2 U3047 ( .A(\PR_add[4][12] ), .B(m1607), .OUT(m2151) );
  XOR2 U3048 ( .A(m2152), .B(m2153), .OUT(N212) );
  XOR2 U3049 ( .A(\PR_add[4][3] ), .B(\PR_mul[6][3] ), .OUT(N211) );
  XOR2 U3050 ( .A(\PR_add[3][19] ), .B(m1619), .OUT(m2154) );
  XOR2 U3051 ( .A(\PR_add[3][18] ), .B(m1620), .OUT(N206) );
  XOR2 U3052 ( .A(m2066), .B(m2065), .OUT(N205) );
  XOR2 U3053 ( .A(\PR_add[3][16] ), .B(m1621), .OUT(m2155) );
  XOR2 U3054 ( .A(m1622), .B(\PR_add[3][15] ), .OUT(N203) );
  XOR2 U3055 ( .A(\PR_add[3][14] ), .B(m1623), .OUT(N202) );
  XOR2 U3056 ( .A(m1625), .B(m1624), .OUT(N201) );
  XOR2 U3057 ( .A(\PR_add[3][12] ), .B(m1626), .OUT(m2156) );
  XOR2 U3058 ( .A(m2157), .B(m2158), .OUT(N189) );
  XOR2 U3059 ( .A(\PR_add[3][0] ), .B(\PR_mul[5][0] ), .OUT(N188) );
  XOR2 U3060 ( .A(\PR_add[2][19] ), .B(m1635), .OUT(N187) );
  XOR2 U3061 ( .A(m1637), .B(m1636), .OUT(N186) );
  XOR2 U3062 ( .A(\PR_add[2][17] ), .B(m1638), .OUT(m2159) );
  XOR2 U3063 ( .A(m1639), .B(\PR_add[2][16] ), .OUT(N184) );
  XOR2 U3064 ( .A(\PR_add[2][15] ), .B(m1640), .OUT(m2160) );
  XOR2 U3065 ( .A(m1641), .B(\PR_add[2][14] ), .OUT(N182) );
  XOR2 U3066 ( .A(\PR_add[2][13] ), .B(m1642), .OUT(N181) );
  XOR2 U3067 ( .A(m1644), .B(m1643), .OUT(N180) );
  XOR2 U3068 ( .A(\PR_add[2][11] ), .B(m1645), .OUT(m2161) );
  XOR2 U3069 ( .A(m2162), .B(m2163), .OUT(N171) );
  XOR2 U3070 ( .A(\PR_add[2][2] ), .B(\PR_mul[4][2] ), .OUT(N170) );
  XOR2 U3071 ( .A(\PR_add[1][19] ), .B(m1656), .OUT(N167) );
  XOR2 U3072 ( .A(m1658), .B(m1657), .OUT(N166) );
  XOR2 U3073 ( .A(\PR_add[1][17] ), .B(m1659), .OUT(m2164) );
  XOR2 U3074 ( .A(m1660), .B(\PR_add[1][16] ), .OUT(N164) );
  XOR2 U3075 ( .A(\PR_add[1][15] ), .B(m2165), .OUT(N163) );
  XOR2 U3076 ( .A(m2077), .B(m2076), .OUT(N162) );
  XOR2 U3077 ( .A(\PR_add[1][13] ), .B(m1661), .OUT(m2166) );
  XOR2 U3078 ( .A(m2169), .B(m2170), .OUT(N129) );
  XOR2 U3079 ( .A(\PR_add[0][0] ), .B(\PR_mul[2][0] ), .OUT(N128) );
  XOR2 U3080 ( .A(m2171), .B(m2172), .OUT(N112) );
  XOR2 U3081 ( .A(\PR_mul[0][3] ), .B(\PR_mul[1][3] ), .OUT(N111) );
  XOR2 U3082 ( .A(\mult_82/ab[1][3] ), .B(m1351), .OUT(m2084) );
  XOR2 U3083 ( .A(m1960), .B(m1961), .OUT(m1696) );
  XOR2 U3084 ( .A(\mult_80/ab[7][0] ), .B(m1379), .OUT(m2086) );
  XOR2 U3085 ( .A(\mult_80/ab[6][0] ), .B(m1971), .OUT(m2087) );
  XOR2 U3086 ( .A(\mult_80/ab[5][0] ), .B(m1965), .OUT(m2088) );
  XOR2 U3087 ( .A(\mult_80/ab[4][0] ), .B(m1373), .OUT(m2089) );
  XOR2 U3088 ( .A(\mult_80/ab[3][0] ), .B(m1962), .OUT(m1697) );
  XOR2 U3089 ( .A(m1369), .B(m1368), .OUT(m2090) );
  XOR2 U3090 ( .A(\mult_76/ab[1][3] ), .B(m1387), .OUT(m2093) );
  XOR2 U3091 ( .A(m1978), .B(m1979), .OUT(m1714) );
  XOR2 U3092 ( .A(\mult_74/ab[7][0] ), .B(m1415), .OUT(m2095) );
  XOR2 U3093 ( .A(\mult_74/ab[6][0] ), .B(m1989), .OUT(m2096) );
  XOR2 U3094 ( .A(\mult_74/ab[5][0] ), .B(m1983), .OUT(m2097) );
  XOR2 U3095 ( .A(\mult_74/ab[4][0] ), .B(m1409), .OUT(m2098) );
  XOR2 U3096 ( .A(\mult_74/ab[3][0] ), .B(m1980), .OUT(m1715) );
  XOR2 U3097 ( .A(m1405), .B(m1404), .OUT(m2099) );
  XOR2 U3098 ( .A(\mult_71/ab[1][3] ), .B(m1423), .OUT(m2102) );
  XOR2 U3099 ( .A(m1996), .B(m1997), .OUT(m1732) );
  XOR2 U3100 ( .A(\mult_69/ab[7][0] ), .B(m1451), .OUT(m2104) );
  XOR2 U3101 ( .A(\mult_69/ab[6][0] ), .B(m2007), .OUT(m2105) );
  XOR2 U3102 ( .A(\mult_69/ab[5][0] ), .B(m2001), .OUT(m2106) );
  XOR2 U3103 ( .A(\mult_69/ab[4][0] ), .B(m1445), .OUT(m2107) );
  XOR2 U3104 ( .A(\mult_69/ab[3][0] ), .B(m1998), .OUT(m1733) );
  XOR2 U3105 ( .A(m1441), .B(m1440), .OUT(m2108) );
  INV U3106 ( .IN(m2071), .OUT(m1639) );
  INV U3107 ( .IN(m2042), .OUT(m1551) );
  INV U3108 ( .IN(m2013), .OUT(m1463) );
  OAI22 U3109 ( .A(m2082), .B(m2173), .C(m1344), .D(m1955), .OUT(m1689) );
  AOI22 U3110 ( .A(\mult_83/ab[2][3] ), .B(\mult_83/ab[3][2] ), .C(m1689), .D(
        m2174), .OUT(m1687) );
  OAI22 U3111 ( .A(m2175), .B(m2176), .C(m1687), .D(m1346), .OUT(m1685) );
  AOI22 U3112 ( .A(\mult_83/ab[4][3] ), .B(\mult_83/ab[5][2] ), .C(m1685), .D(
        m2177), .OUT(m1683) );
  OAI22 U3113 ( .A(m2178), .B(m2179), .C(m1683), .D(m1348), .OUT(m1681) );
  AOI22 U3114 ( .A(\mult_83/ab[6][3] ), .B(\mult_83/ab[7][2] ), .C(m1681), .D(
        m2180), .OUT(m1338) );
  AOI22 U3115 ( .A(m2181), .B(\mult_82/ab[7][0] ), .C(m1358), .D(
        \mult_82/ab[4][3] ), .OUT(m1316) );
  OAI22 U3116 ( .A(m1695), .B(m1961), .C(m1361), .D(m1960), .OUT(m2182) );
  AOI22 U3117 ( .A(\mult_80/ab[2][2] ), .B(\mult_80/ab[3][1] ), .C(m2182), .D(
        m2184), .OUT(m2183) );
  OAI22 U3118 ( .A(m2186), .B(m2187), .C(m2183), .D(m1363), .OUT(m2185) );
  AOI22 U3119 ( .A(\mult_80/ab[4][2] ), .B(\mult_80/ab[5][1] ), .C(m2185), .D(
        m2189), .OUT(m2188) );
  OAI22 U3120 ( .A(m2191), .B(m2192), .C(m2188), .D(m1365), .OUT(m2190) );
  AOI22 U3121 ( .A(\mult_80/ab[6][2] ), .B(\mult_80/ab[7][1] ), .C(m2190), .D(
        m2193), .OUT(m1334) );
  INV U3122 ( .IN(m1377), .OUT(m1971) );
  AOI22 U3123 ( .A(m1379), .B(\mult_80/ab[7][0] ), .C(m2194), .D(m2085), .OUT(
        m1336) );
  OAI22 U3124 ( .A(m2091), .B(m2195), .C(m1380), .D(m1973), .OUT(m1707) );
  AOI22 U3125 ( .A(\mult_77/ab[2][3] ), .B(\mult_77/ab[3][2] ), .C(m1707), .D(
        m2196), .OUT(m1705) );
  OAI22 U3126 ( .A(m2197), .B(m2198), .C(m1705), .D(m1382), .OUT(m1703) );
  AOI22 U3127 ( .A(\mult_77/ab[4][3] ), .B(\mult_77/ab[5][2] ), .C(m1703), .D(
        m2199), .OUT(m1701) );
  OAI22 U3128 ( .A(m2200), .B(m2201), .C(m1701), .D(m1384), .OUT(m1699) );
  AOI22 U3129 ( .A(\mult_77/ab[6][3] ), .B(\mult_77/ab[7][2] ), .C(m1699), .D(
        m2202), .OUT(m1332) );
  AOI22 U3130 ( .A(m2203), .B(\mult_76/ab[7][0] ), .C(m1394), .D(
        \mult_76/ab[4][3] ), .OUT(m1330) );
  OAI22 U3131 ( .A(m1713), .B(m1979), .C(m1397), .D(m1978), .OUT(m2204) );
  AOI22 U3132 ( .A(\mult_74/ab[2][2] ), .B(\mult_74/ab[3][1] ), .C(m2204), .D(
        m2206), .OUT(m2205) );
  OAI22 U3133 ( .A(m2208), .B(m2209), .C(m2205), .D(m1399), .OUT(m2207) );
  AOI22 U3134 ( .A(\mult_74/ab[4][2] ), .B(\mult_74/ab[5][1] ), .C(m2207), .D(
        m2211), .OUT(m2210) );
  OAI22 U3135 ( .A(m2213), .B(m2214), .C(m2210), .D(m1401), .OUT(m2212) );
  AOI22 U3136 ( .A(\mult_74/ab[6][2] ), .B(\mult_74/ab[7][1] ), .C(m2212), .D(
        m2215), .OUT(m1326) );
  INV U3137 ( .IN(m1413), .OUT(m1989) );
  AOI22 U3138 ( .A(m1415), .B(\mult_74/ab[7][0] ), .C(m2216), .D(m2094), .OUT(
        m1328) );
  OAI22 U3139 ( .A(m2100), .B(m2217), .C(m1416), .D(m1991), .OUT(m1725) );
  AOI22 U3140 ( .A(\mult_72/ab[2][3] ), .B(\mult_72/ab[3][2] ), .C(m1725), .D(
        m2218), .OUT(m1723) );
  OAI22 U3141 ( .A(m2219), .B(m2220), .C(m1723), .D(m1418), .OUT(m1721) );
  AOI22 U3142 ( .A(\mult_72/ab[4][3] ), .B(\mult_72/ab[5][2] ), .C(m1721), .D(
        m2221), .OUT(m1719) );
  OAI22 U3143 ( .A(m2222), .B(m2223), .C(m1719), .D(m1420), .OUT(m1717) );
  AOI22 U3144 ( .A(\mult_72/ab[6][3] ), .B(\mult_72/ab[7][2] ), .C(m1717), .D(
        m2224), .OUT(m1324) );
  AOI22 U3145 ( .A(m2225), .B(\mult_71/ab[7][0] ), .C(m1430), .D(
        \mult_71/ab[4][3] ), .OUT(m1322) );
  OAI22 U3146 ( .A(m1731), .B(m1997), .C(m1433), .D(m1996), .OUT(m2226) );
  AOI22 U3147 ( .A(\mult_69/ab[2][2] ), .B(\mult_69/ab[3][1] ), .C(m2226), .D(
        m2228), .OUT(m2227) );
  OAI22 U3148 ( .A(m2230), .B(m2231), .C(m2227), .D(m1435), .OUT(m2229) );
  AOI22 U3149 ( .A(\mult_69/ab[4][2] ), .B(\mult_69/ab[5][1] ), .C(m2229), .D(
        m2233), .OUT(m2232) );
  OAI22 U3150 ( .A(m2235), .B(m2236), .C(m2232), .D(m1437), .OUT(m2234) );
  AOI22 U3151 ( .A(\mult_69/ab[6][2] ), .B(\mult_69/ab[7][1] ), .C(m2234), .D(
        m2237), .OUT(m1318) );
  INV U3152 ( .IN(m1449), .OUT(m2007) );
  AOI22 U3153 ( .A(m1451), .B(\mult_69/ab[7][0] ), .C(m2238), .D(m2103), .OUT(
        m1320) );
  OAI22 U3154 ( .A(m2112), .B(m2239), .C(m1452), .D(m2009), .OUT(m1745) );
  AOI22 U3155 ( .A(\PR_mul[14][4] ), .B(\PR_add[12][4] ), .C(m1745), .D(m2240), 
        .OUT(m1743) );
  OAI22 U3156 ( .A(m2241), .B(m2242), .C(m1743), .D(m1454), .OUT(m1741) );
  AOI22 U3157 ( .A(\PR_mul[14][6] ), .B(\PR_add[12][6] ), .C(m1741), .D(m2243), 
        .OUT(m1739) );
  OAI22 U3158 ( .A(m2244), .B(m2245), .C(m1739), .D(m1456), .OUT(m1737) );
  AOI22 U3159 ( .A(\PR_mul[14][8] ), .B(\PR_add[12][8] ), .C(m1737), .D(m2246), 
        .OUT(m1735) );
  OAI22 U3160 ( .A(m2010), .B(m2011), .C(m1735), .D(m1458), .OUT(m1470) );
  OAI22 U3161 ( .A(m2247), .B(m2248), .C(m1763), .D(m1471), .OUT(m1761) );
  AOI22 U3162 ( .A(\PR_mul[13][4] ), .B(\PR_add[11][4] ), .C(m1761), .D(m2249), 
        .OUT(m1759) );
  OAI22 U3163 ( .A(m2250), .B(m2251), .C(m1759), .D(m1473), .OUT(m1757) );
  AOI22 U3164 ( .A(\PR_mul[13][6] ), .B(\PR_add[11][6] ), .C(m1757), .D(m2252), 
        .OUT(m1755) );
  OAI22 U3165 ( .A(m2253), .B(m2254), .C(m1755), .D(m1475), .OUT(m1753) );
  AOI22 U3166 ( .A(\PR_mul[13][8] ), .B(\PR_add[11][8] ), .C(m1753), .D(m2255), 
        .OUT(m1751) );
  OAI22 U3167 ( .A(m2256), .B(m2257), .C(m1751), .D(m1477), .OUT(m1749) );
  AOI22 U3168 ( .A(\PR_mul[13][10] ), .B(\PR_add[11][10] ), .C(m1749), .D(
        m2258), .OUT(m1747) );
  OAI22 U3169 ( .A(m2015), .B(m2016), .C(m1747), .D(m1479), .OUT(m1486) );
  NOR2 U3170 ( .A(m2019), .B(m2018), .OUT(m2115) );
  OAI22 U3171 ( .A(m2122), .B(m2259), .C(m1487), .D(m2020), .OUT(m1783) );
  AOI22 U3172 ( .A(\PR_mul[12][2] ), .B(\PR_add[10][2] ), .C(m1783), .D(m2260), 
        .OUT(m1781) );
  OAI22 U3173 ( .A(m2261), .B(m2262), .C(m1781), .D(m1489), .OUT(m1779) );
  AOI22 U3174 ( .A(\PR_mul[12][4] ), .B(\PR_add[10][4] ), .C(m1779), .D(m2263), 
        .OUT(m1777) );
  OAI22 U3175 ( .A(m2264), .B(m2265), .C(m1777), .D(m1491), .OUT(m1775) );
  AOI22 U3176 ( .A(\PR_mul[12][6] ), .B(\PR_add[10][6] ), .C(m1775), .D(m2266), 
        .OUT(m1773) );
  OAI22 U3177 ( .A(m2267), .B(m2268), .C(m1773), .D(m1493), .OUT(m1771) );
  AOI22 U3178 ( .A(\PR_mul[12][8] ), .B(\PR_add[10][8] ), .C(m1771), .D(m2269), 
        .OUT(m1769) );
  OAI22 U3179 ( .A(m2270), .B(m2271), .C(m1769), .D(m1495), .OUT(m1767) );
  AOI22 U3180 ( .A(\PR_mul[12][10] ), .B(\PR_add[10][10] ), .C(m1767), .D(
        m2272), .OUT(m1765) );
  OAI22 U3181 ( .A(m2021), .B(m2022), .C(m1765), .D(m1497), .OUT(m1504) );
  NOR2 U3182 ( .A(m2025), .B(m2024), .OUT(m2120) );
  OAI22 U3183 ( .A(m2127), .B(m2273), .C(m1505), .D(m2026), .OUT(m1795) );
  AOI22 U3184 ( .A(\PR_mul[11][5] ), .B(\PR_add[9][5] ), .C(m1795), .D(m2274), 
        .OUT(m1793) );
  OAI22 U3185 ( .A(m2275), .B(m2276), .C(m1793), .D(m1507), .OUT(m1791) );
  AOI22 U3186 ( .A(\PR_mul[11][7] ), .B(\PR_add[9][7] ), .C(m1791), .D(m2277), 
        .OUT(m1789) );
  OAI22 U3187 ( .A(m2278), .B(m2279), .C(m1789), .D(m1509), .OUT(m1787) );
  AOI22 U3188 ( .A(\PR_mul[11][9] ), .B(\PR_add[9][9] ), .C(m1787), .D(m2280), 
        .OUT(m1785) );
  OAI22 U3189 ( .A(m2027), .B(m2028), .C(m1785), .D(m1511), .OUT(m1520) );
  OAI22 U3190 ( .A(m2132), .B(m2281), .C(m1521), .D(m2032), .OUT(m1813) );
  AOI22 U3191 ( .A(\PR_mul[10][2] ), .B(\PR_add[8][2] ), .C(m1813), .D(m2282), 
        .OUT(m1811) );
  OAI22 U3192 ( .A(m2283), .B(m2284), .C(m1811), .D(m1523), .OUT(m1809) );
  AOI22 U3193 ( .A(\PR_mul[10][4] ), .B(\PR_add[8][4] ), .C(m1809), .D(m2285), 
        .OUT(m1807) );
  OAI22 U3194 ( .A(m2286), .B(m2287), .C(m1807), .D(m1525), .OUT(m1805) );
  AOI22 U3195 ( .A(\PR_mul[10][6] ), .B(\PR_add[8][6] ), .C(m1805), .D(m2288), 
        .OUT(m1803) );
  OAI22 U3196 ( .A(m2289), .B(m2290), .C(m1803), .D(m1527), .OUT(m1801) );
  AOI22 U3197 ( .A(\PR_mul[10][8] ), .B(\PR_add[8][8] ), .C(m1801), .D(m2292), 
        .OUT(m2291) );
  AOI22 U3198 ( .A(\PR_mul[10][9] ), .B(\PR_add[8][9] ), .C(m1799), .D(m2293), 
        .OUT(m1797) );
  OAI22 U3199 ( .A(m2033), .B(m2034), .C(m1797), .D(m1530), .OUT(m1539) );
  OAI22 U3200 ( .A(m2137), .B(m2294), .C(m1540), .D(m2038), .OUT(m1825) );
  AOI22 U3201 ( .A(\PR_mul[9][4] ), .B(\PR_add[7][4] ), .C(m1825), .D(m2295), 
        .OUT(m1823) );
  OAI22 U3202 ( .A(m2296), .B(m2297), .C(m1823), .D(m1542), .OUT(m1821) );
  AOI22 U3203 ( .A(\PR_mul[9][6] ), .B(\PR_add[7][6] ), .C(m1821), .D(m2298), 
        .OUT(m1819) );
  OAI22 U3204 ( .A(m2299), .B(m2300), .C(m1819), .D(m1544), .OUT(m1817) );
  AOI22 U3205 ( .A(\PR_mul[9][8] ), .B(\PR_add[7][8] ), .C(m1817), .D(m2301), 
        .OUT(m1815) );
  OAI22 U3206 ( .A(m2039), .B(m2040), .C(m1815), .D(m1546), .OUT(m1558) );
  OAI22 U3207 ( .A(m2302), .B(m2303), .C(m1843), .D(m1559), .OUT(m1841) );
  AOI22 U3208 ( .A(\PR_mul[8][4] ), .B(\PR_add[6][4] ), .C(m1841), .D(m2304), 
        .OUT(m1839) );
  OAI22 U3209 ( .A(m2305), .B(m2306), .C(m1839), .D(m1561), .OUT(m1837) );
  AOI22 U3210 ( .A(\PR_mul[8][6] ), .B(\PR_add[6][6] ), .C(m1837), .D(m2307), 
        .OUT(m1835) );
  OAI22 U3211 ( .A(m2308), .B(m2309), .C(m1835), .D(m1563), .OUT(m1833) );
  AOI22 U3212 ( .A(\PR_mul[8][8] ), .B(\PR_add[6][8] ), .C(m1833), .D(m2310), 
        .OUT(m1831) );
  OAI22 U3213 ( .A(m2311), .B(m2312), .C(m1831), .D(m1565), .OUT(m1829) );
  AOI22 U3214 ( .A(\PR_mul[8][10] ), .B(\PR_add[6][10] ), .C(m1829), .D(m2313), 
        .OUT(m1827) );
  OAI22 U3215 ( .A(m2044), .B(m2045), .C(m1827), .D(m1567), .OUT(m1574) );
  NOR2 U3216 ( .A(m2048), .B(m2047), .OUT(m2140) );
  OAI22 U3217 ( .A(m2147), .B(m2314), .C(m1575), .D(m2049), .OUT(m1863) );
  AOI22 U3218 ( .A(\PR_mul[7][2] ), .B(\PR_add[5][2] ), .C(m1863), .D(m2315), 
        .OUT(m1861) );
  OAI22 U3219 ( .A(m2316), .B(m2317), .C(m1861), .D(m1577), .OUT(m1859) );
  AOI22 U3220 ( .A(\PR_mul[7][4] ), .B(\PR_add[5][4] ), .C(m1859), .D(m2318), 
        .OUT(m1857) );
  OAI22 U3221 ( .A(m2319), .B(m2320), .C(m1857), .D(m1579), .OUT(m1855) );
  AOI22 U3222 ( .A(\PR_mul[7][6] ), .B(\PR_add[5][6] ), .C(m1855), .D(m2321), 
        .OUT(m1853) );
  OAI22 U3223 ( .A(m2322), .B(m2323), .C(m1853), .D(m1581), .OUT(m1851) );
  AOI22 U3224 ( .A(\PR_mul[7][8] ), .B(\PR_add[5][8] ), .C(m1851), .D(m2324), 
        .OUT(m1849) );
  OAI22 U3225 ( .A(m2325), .B(m2326), .C(m1849), .D(m1583), .OUT(m1847) );
  AOI22 U3226 ( .A(\PR_mul[7][10] ), .B(\PR_add[5][10] ), .C(m1847), .D(m2327), 
        .OUT(m1845) );
  OAI22 U3227 ( .A(m2050), .B(m2051), .C(m1845), .D(m1585), .OUT(m1592) );
  NOR2 U3228 ( .A(m2054), .B(m2053), .OUT(m2145) );
  OAI22 U3229 ( .A(m2152), .B(m2328), .C(m1593), .D(m2055), .OUT(m1875) );
  AOI22 U3230 ( .A(\PR_mul[6][5] ), .B(\PR_add[4][5] ), .C(m1875), .D(m2329), 
        .OUT(m1873) );
  OAI22 U3231 ( .A(m2330), .B(m2331), .C(m1873), .D(m1595), .OUT(m1871) );
  AOI22 U3232 ( .A(\PR_mul[6][7] ), .B(\PR_add[4][7] ), .C(m1871), .D(m2332), 
        .OUT(m1869) );
  OAI22 U3233 ( .A(m2333), .B(m2334), .C(m1869), .D(m1597), .OUT(m1867) );
  AOI22 U3234 ( .A(\PR_mul[6][9] ), .B(\PR_add[4][9] ), .C(m1867), .D(m2335), 
        .OUT(m1865) );
  OAI22 U3235 ( .A(m2056), .B(m2057), .C(m1865), .D(m1599), .OUT(m1608) );
  OAI22 U3236 ( .A(m2157), .B(m2336), .C(m1609), .D(m2061), .OUT(m1893) );
  AOI22 U3237 ( .A(\PR_mul[5][2] ), .B(\PR_add[3][2] ), .C(m1893), .D(m2337), 
        .OUT(m1891) );
  OAI22 U3238 ( .A(m2338), .B(m2339), .C(m1891), .D(m1611), .OUT(m1889) );
  AOI22 U3239 ( .A(\PR_mul[5][4] ), .B(\PR_add[3][4] ), .C(m1889), .D(m2340), 
        .OUT(m1887) );
  OAI22 U3240 ( .A(m2341), .B(m2342), .C(m1887), .D(m1613), .OUT(m1885) );
  AOI22 U3241 ( .A(\PR_mul[5][6] ), .B(\PR_add[3][6] ), .C(m1885), .D(m2343), 
        .OUT(m1883) );
  OAI22 U3242 ( .A(m2344), .B(m2345), .C(m1883), .D(m1615), .OUT(m1881) );
  AOI22 U3243 ( .A(\PR_mul[5][8] ), .B(\PR_add[3][8] ), .C(m1881), .D(m2347), 
        .OUT(m2346) );
  AOI22 U3244 ( .A(\PR_mul[5][9] ), .B(\PR_add[3][9] ), .C(m1879), .D(m2348), 
        .OUT(m1877) );
  OAI22 U3245 ( .A(m2062), .B(m2063), .C(m1877), .D(m1618), .OUT(m1627) );
  OAI22 U3246 ( .A(m2162), .B(m2349), .C(m1628), .D(m2067), .OUT(m1905) );
  AOI22 U3247 ( .A(\PR_mul[4][4] ), .B(\PR_add[2][4] ), .C(m1905), .D(m2350), 
        .OUT(m1903) );
  OAI22 U3248 ( .A(m2351), .B(m2352), .C(m1903), .D(m1630), .OUT(m1901) );
  AOI22 U3249 ( .A(\PR_mul[4][6] ), .B(\PR_add[2][6] ), .C(m1901), .D(m2353), 
        .OUT(m1899) );
  OAI22 U3250 ( .A(m2354), .B(m2355), .C(m1899), .D(m1632), .OUT(m1897) );
  AOI22 U3251 ( .A(\PR_mul[4][8] ), .B(\PR_add[2][8] ), .C(m1897), .D(m2356), 
        .OUT(m1895) );
  OAI22 U3252 ( .A(m2068), .B(m2069), .C(m1895), .D(m1634), .OUT(m1646) );
  OAI22 U3253 ( .A(m2357), .B(m2358), .C(m1923), .D(m1647), .OUT(m1921) );
  AOI22 U3254 ( .A(\PR_mul[3][4] ), .B(\PR_add[1][4] ), .C(m1921), .D(m2359), 
        .OUT(m1919) );
  OAI22 U3255 ( .A(m2360), .B(m2361), .C(m1919), .D(m1649), .OUT(m1917) );
  AOI22 U3256 ( .A(\PR_mul[3][6] ), .B(\PR_add[1][6] ), .C(m1917), .D(m2362), 
        .OUT(m1915) );
  OAI22 U3257 ( .A(m2363), .B(m2364), .C(m1915), .D(m1651), .OUT(m1913) );
  AOI22 U3258 ( .A(\PR_mul[3][8] ), .B(\PR_add[1][8] ), .C(m1913), .D(m2365), 
        .OUT(m1911) );
  OAI22 U3259 ( .A(m2366), .B(m2367), .C(m1911), .D(m1653), .OUT(m1909) );
  AOI22 U3260 ( .A(\PR_mul[3][10] ), .B(\PR_add[1][10] ), .C(m1909), .D(m2368), 
        .OUT(m1907) );
  OAI22 U3261 ( .A(m2073), .B(m2074), .C(m1907), .D(m1655), .OUT(m1662) );
  NOR2 U3262 ( .A(m2077), .B(m2076), .OUT(m2165) );
  OAI22 U3263 ( .A(m2169), .B(m2369), .C(m1663), .D(m2078), .OUT(m1943) );
  AOI22 U3264 ( .A(\PR_mul[2][2] ), .B(\PR_add[0][2] ), .C(m1943), .D(m2370), 
        .OUT(m1941) );
  OAI22 U3265 ( .A(m2371), .B(m2372), .C(m1941), .D(m1665), .OUT(m1939) );
  AOI22 U3266 ( .A(\PR_mul[2][4] ), .B(\PR_add[0][4] ), .C(m1939), .D(m2373), 
        .OUT(m1937) );
  OAI22 U3267 ( .A(m2374), .B(m2375), .C(m1937), .D(m1667), .OUT(m1935) );
  AOI22 U3268 ( .A(\PR_mul[2][6] ), .B(\PR_add[0][6] ), .C(m1935), .D(m2376), 
        .OUT(m1933) );
  OAI22 U3269 ( .A(m2377), .B(m2378), .C(m1933), .D(m1669), .OUT(m1931) );
  AOI22 U3270 ( .A(\PR_mul[2][8] ), .B(\PR_add[0][8] ), .C(m1931), .D(m2379), 
        .OUT(m1929) );
  OAI22 U3271 ( .A(m2380), .B(m2381), .C(m1929), .D(m1671), .OUT(m1927) );
  AOI22 U3272 ( .A(\PR_mul[2][10] ), .B(\PR_add[0][10] ), .C(m1927), .D(m2382), 
        .OUT(m1925) );
  OAI22 U3273 ( .A(m2079), .B(m2080), .C(m1925), .D(m1673), .OUT(N140) );
  OAI22 U3274 ( .A(m2171), .B(m2383), .C(m1674), .D(m2081), .OUT(m1954) );
  AOI22 U3275 ( .A(\PR_mul[1][5] ), .B(\PR_mul[0][5] ), .C(m1954), .D(m2384), 
        .OUT(m1952) );
  OAI22 U3276 ( .A(m2385), .B(m2386), .C(m1952), .D(m1676), .OUT(m1950) );
  AOI22 U3277 ( .A(\PR_mul[1][7] ), .B(\PR_mul[0][7] ), .C(m1950), .D(m2387), 
        .OUT(m1948) );
  OAI22 U3278 ( .A(m2388), .B(m2389), .C(m1948), .D(m1678), .OUT(m1946) );
  AOI22 U3279 ( .A(\PR_mul[1][9] ), .B(\PR_mul[0][9] ), .C(m1946), .D(m2390), 
        .OUT(m1342) );
  XOR2 U3280 ( .A(m2391), .B(m2182), .OUT(m1967) );
  XOR2 U3281 ( .A(m2392), .B(m2183), .OUT(m1969) );
  XOR2 U3282 ( .A(m2394), .B(m2185), .OUT(m2393) );
  XOR2 U3283 ( .A(m2395), .B(m2188), .OUT(m2085) );
  XOR2 U3284 ( .A(m2397), .B(m2190), .OUT(m2396) );
  XOR2 U3285 ( .A(m2398), .B(m2204), .OUT(m1985) );
  XOR2 U3286 ( .A(m2399), .B(m2205), .OUT(m1987) );
  XOR2 U3287 ( .A(m2401), .B(m2207), .OUT(m2400) );
  XOR2 U3288 ( .A(m2402), .B(m2210), .OUT(m2094) );
  XOR2 U3289 ( .A(m2404), .B(m2212), .OUT(m2403) );
  XOR2 U3290 ( .A(m2405), .B(m2226), .OUT(m2003) );
  XOR2 U3291 ( .A(m2406), .B(m2227), .OUT(m2005) );
  XOR2 U3292 ( .A(m2408), .B(m2229), .OUT(m2407) );
  XOR2 U3293 ( .A(m2409), .B(m2232), .OUT(m2103) );
  XOR2 U3294 ( .A(m2411), .B(m2234), .OUT(m2410) );
  XOR2 U3295 ( .A(\mult_83/ab[6][3] ), .B(\mult_83/ab[7][2] ), .OUT(m1680) );
  XOR2 U3296 ( .A(m2178), .B(\mult_83/ab[6][2] ), .OUT(m1682) );
  XOR2 U3297 ( .A(\mult_83/ab[4][3] ), .B(\mult_83/ab[5][2] ), .OUT(m1684) );
  XOR2 U3298 ( .A(m2175), .B(\mult_83/ab[4][2] ), .OUT(m1686) );
  XOR2 U3299 ( .A(\mult_83/ab[2][3] ), .B(\mult_83/ab[3][2] ), .OUT(m1688) );
  XOR2 U3300 ( .A(m1955), .B(\mult_83/ab[2][2] ), .OUT(m2083) );
  XOR2 U3301 ( .A(m1359), .B(\mult_82/ab[4][3] ), .OUT(m1690) );
  XOR2 U3302 ( .A(m1356), .B(\mult_82/ab[3][3] ), .OUT(m1691) );
  XOR2 U3303 ( .A(m1353), .B(\mult_82/ab[2][3] ), .OUT(m1692) );
  XOR2 U3304 ( .A(\mult_80/ab[2][2] ), .B(\mult_80/ab[3][1] ), .OUT(m2391) );
  XOR2 U3305 ( .A(m2186), .B(m2187), .OUT(m2392) );
  XOR2 U3306 ( .A(\mult_80/ab[4][2] ), .B(\mult_80/ab[5][1] ), .OUT(m2394) );
  XOR2 U3307 ( .A(m2191), .B(\mult_80/ab[6][1] ), .OUT(m2395) );
  XOR2 U3308 ( .A(\mult_80/ab[6][2] ), .B(\mult_80/ab[7][1] ), .OUT(m2397) );
  XOR2 U3309 ( .A(\mult_77/ab[6][3] ), .B(\mult_77/ab[7][2] ), .OUT(m1698) );
  XOR2 U3310 ( .A(m2200), .B(\mult_77/ab[6][2] ), .OUT(m1700) );
  XOR2 U3311 ( .A(\mult_77/ab[4][3] ), .B(\mult_77/ab[5][2] ), .OUT(m1702) );
  XOR2 U3312 ( .A(m2197), .B(\mult_77/ab[4][2] ), .OUT(m1704) );
  XOR2 U3313 ( .A(\mult_77/ab[2][3] ), .B(\mult_77/ab[3][2] ), .OUT(m1706) );
  XOR2 U3314 ( .A(m1973), .B(\mult_77/ab[2][2] ), .OUT(m2092) );
  XOR2 U3315 ( .A(m1395), .B(\mult_76/ab[4][3] ), .OUT(m1708) );
  XOR2 U3316 ( .A(m1392), .B(\mult_76/ab[3][3] ), .OUT(m1709) );
  XOR2 U3317 ( .A(m1389), .B(\mult_76/ab[2][3] ), .OUT(m1710) );
  XOR2 U3318 ( .A(\mult_74/ab[2][2] ), .B(\mult_74/ab[3][1] ), .OUT(m2398) );
  XOR2 U3319 ( .A(m2208), .B(m2209), .OUT(m2399) );
  XOR2 U3320 ( .A(\mult_74/ab[4][2] ), .B(\mult_74/ab[5][1] ), .OUT(m2401) );
  XOR2 U3321 ( .A(m2213), .B(\mult_74/ab[6][1] ), .OUT(m2402) );
  XOR2 U3322 ( .A(\mult_74/ab[6][2] ), .B(\mult_74/ab[7][1] ), .OUT(m2404) );
  XOR2 U3323 ( .A(\mult_72/ab[6][3] ), .B(\mult_72/ab[7][2] ), .OUT(m1716) );
  XOR2 U3324 ( .A(m2222), .B(\mult_72/ab[6][2] ), .OUT(m1718) );
  XOR2 U3325 ( .A(\mult_72/ab[4][3] ), .B(\mult_72/ab[5][2] ), .OUT(m1720) );
  XOR2 U3326 ( .A(m2219), .B(\mult_72/ab[4][2] ), .OUT(m1722) );
  XOR2 U3327 ( .A(\mult_72/ab[2][3] ), .B(\mult_72/ab[3][2] ), .OUT(m1724) );
  XOR2 U3328 ( .A(m1991), .B(\mult_72/ab[2][2] ), .OUT(m2101) );
  XOR2 U3329 ( .A(m1431), .B(\mult_71/ab[4][3] ), .OUT(m1726) );
  XOR2 U3330 ( .A(m1428), .B(\mult_71/ab[3][3] ), .OUT(m1727) );
  XOR2 U3331 ( .A(m1425), .B(\mult_71/ab[2][3] ), .OUT(m1728) );
  XOR2 U3332 ( .A(\mult_69/ab[2][2] ), .B(\mult_69/ab[3][1] ), .OUT(m2405) );
  XOR2 U3333 ( .A(m2230), .B(m2231), .OUT(m2406) );
  XOR2 U3334 ( .A(\mult_69/ab[4][2] ), .B(\mult_69/ab[5][1] ), .OUT(m2408) );
  XOR2 U3335 ( .A(m2235), .B(\mult_69/ab[6][1] ), .OUT(m2409) );
  XOR2 U3336 ( .A(\mult_69/ab[6][2] ), .B(\mult_69/ab[7][1] ), .OUT(m2411) );
  XOR2 U3337 ( .A(m2010), .B(\PR_add[12][9] ), .OUT(m1734) );
  XOR2 U3338 ( .A(\PR_mul[14][8] ), .B(\PR_add[12][8] ), .OUT(m1736) );
  XOR2 U3339 ( .A(m2244), .B(\PR_add[12][7] ), .OUT(m1738) );
  XOR2 U3340 ( .A(\PR_mul[14][6] ), .B(\PR_add[12][6] ), .OUT(m1740) );
  XOR2 U3341 ( .A(m2241), .B(\PR_add[12][5] ), .OUT(m1742) );
  XOR2 U3342 ( .A(\PR_mul[14][4] ), .B(\PR_add[12][4] ), .OUT(m1744) );
  XOR2 U3343 ( .A(m2009), .B(\PR_add[12][3] ), .OUT(m2113) );
  XOR2 U3344 ( .A(m2015), .B(\PR_add[11][11] ), .OUT(m1746) );
  XOR2 U3345 ( .A(\PR_mul[13][10] ), .B(\PR_add[11][10] ), .OUT(m1748) );
  XOR2 U3346 ( .A(m2256), .B(\PR_add[11][9] ), .OUT(m1750) );
  XOR2 U3347 ( .A(\PR_mul[13][8] ), .B(\PR_add[11][8] ), .OUT(m1752) );
  XOR2 U3348 ( .A(m2253), .B(\PR_add[11][7] ), .OUT(m1754) );
  XOR2 U3349 ( .A(\PR_mul[13][6] ), .B(\PR_add[11][6] ), .OUT(m1756) );
  XOR2 U3350 ( .A(m2250), .B(\PR_add[11][5] ), .OUT(m1758) );
  XOR2 U3351 ( .A(\PR_mul[13][4] ), .B(\PR_add[11][4] ), .OUT(m1760) );
  XOR2 U3352 ( .A(m2247), .B(\PR_add[11][3] ), .OUT(m1762) );
  XOR2 U3353 ( .A(\PR_mul[13][2] ), .B(\PR_add[11][2] ), .OUT(N350) );
  XOR2 U3354 ( .A(m2021), .B(\PR_add[10][11] ), .OUT(m1764) );
  XOR2 U3355 ( .A(\PR_mul[12][10] ), .B(\PR_add[10][10] ), .OUT(m1766) );
  XOR2 U3356 ( .A(m2270), .B(\PR_add[10][9] ), .OUT(m1768) );
  XOR2 U3357 ( .A(\PR_mul[12][8] ), .B(\PR_add[10][8] ), .OUT(m1770) );
  XOR2 U3358 ( .A(m2267), .B(\PR_add[10][7] ), .OUT(m1772) );
  XOR2 U3359 ( .A(\PR_mul[12][6] ), .B(\PR_add[10][6] ), .OUT(m1774) );
  XOR2 U3360 ( .A(m2264), .B(\PR_add[10][5] ), .OUT(m1776) );
  XOR2 U3361 ( .A(\PR_mul[12][4] ), .B(\PR_add[10][4] ), .OUT(m1778) );
  XOR2 U3362 ( .A(m2261), .B(\PR_add[10][3] ), .OUT(m1780) );
  XOR2 U3363 ( .A(\PR_mul[12][2] ), .B(\PR_add[10][2] ), .OUT(m1782) );
  XOR2 U3364 ( .A(m2020), .B(\PR_add[10][1] ), .OUT(m2123) );
  XOR2 U3365 ( .A(m2027), .B(\PR_add[9][10] ), .OUT(m1784) );
  XOR2 U3366 ( .A(\PR_mul[11][9] ), .B(\PR_add[9][9] ), .OUT(m1786) );
  XOR2 U3367 ( .A(m2278), .B(\PR_add[9][8] ), .OUT(m1788) );
  XOR2 U3368 ( .A(\PR_mul[11][7] ), .B(\PR_add[9][7] ), .OUT(m1790) );
  XOR2 U3369 ( .A(m2275), .B(\PR_add[9][6] ), .OUT(m1792) );
  XOR2 U3370 ( .A(\PR_mul[11][5] ), .B(\PR_add[9][5] ), .OUT(m1794) );
  XOR2 U3371 ( .A(m2026), .B(\PR_add[9][4] ), .OUT(m2128) );
  XOR2 U3372 ( .A(m2033), .B(\PR_add[8][10] ), .OUT(m1796) );
  XOR2 U3373 ( .A(\PR_mul[10][9] ), .B(\PR_add[8][9] ), .OUT(m1798) );
  XOR2 U3374 ( .A(\PR_mul[10][8] ), .B(\PR_add[8][8] ), .OUT(m1800) );
  XOR2 U3375 ( .A(m2289), .B(\PR_add[8][7] ), .OUT(m1802) );
  XOR2 U3376 ( .A(\PR_mul[10][6] ), .B(\PR_add[8][6] ), .OUT(m1804) );
  XOR2 U3377 ( .A(m2286), .B(\PR_add[8][5] ), .OUT(m1806) );
  XOR2 U3378 ( .A(\PR_mul[10][4] ), .B(\PR_add[8][4] ), .OUT(m1808) );
  XOR2 U3379 ( .A(m2283), .B(\PR_add[8][3] ), .OUT(m1810) );
  XOR2 U3380 ( .A(\PR_mul[10][2] ), .B(\PR_add[8][2] ), .OUT(m1812) );
  XOR2 U3381 ( .A(m2032), .B(\PR_add[8][1] ), .OUT(m2133) );
  XOR2 U3382 ( .A(m2039), .B(\PR_add[7][9] ), .OUT(m1814) );
  XOR2 U3383 ( .A(\PR_mul[9][8] ), .B(\PR_add[7][8] ), .OUT(m1816) );
  XOR2 U3384 ( .A(m2299), .B(\PR_add[7][7] ), .OUT(m1818) );
  XOR2 U3385 ( .A(\PR_mul[9][6] ), .B(\PR_add[7][6] ), .OUT(m1820) );
  XOR2 U3386 ( .A(m2296), .B(\PR_add[7][5] ), .OUT(m1822) );
  XOR2 U3387 ( .A(\PR_mul[9][4] ), .B(\PR_add[7][4] ), .OUT(m1824) );
  XOR2 U3388 ( .A(m2038), .B(\PR_add[7][3] ), .OUT(m2138) );
  XOR2 U3389 ( .A(m2044), .B(\PR_add[6][11] ), .OUT(m1826) );
  XOR2 U3390 ( .A(\PR_mul[8][10] ), .B(\PR_add[6][10] ), .OUT(m1828) );
  XOR2 U3391 ( .A(m2311), .B(\PR_add[6][9] ), .OUT(m1830) );
  XOR2 U3392 ( .A(\PR_mul[8][8] ), .B(\PR_add[6][8] ), .OUT(m1832) );
  XOR2 U3393 ( .A(m2308), .B(\PR_add[6][7] ), .OUT(m1834) );
  XOR2 U3394 ( .A(\PR_mul[8][6] ), .B(\PR_add[6][6] ), .OUT(m1836) );
  XOR2 U3395 ( .A(m2305), .B(\PR_add[6][5] ), .OUT(m1838) );
  XOR2 U3396 ( .A(\PR_mul[8][4] ), .B(\PR_add[6][4] ), .OUT(m1840) );
  XOR2 U3397 ( .A(m2302), .B(\PR_add[6][3] ), .OUT(m1842) );
  XOR2 U3398 ( .A(\PR_mul[8][2] ), .B(\PR_add[6][2] ), .OUT(N250) );
  XOR2 U3399 ( .A(m2050), .B(\PR_add[5][11] ), .OUT(m1844) );
  XOR2 U3400 ( .A(\PR_mul[7][10] ), .B(\PR_add[5][10] ), .OUT(m1846) );
  XOR2 U3401 ( .A(m2325), .B(\PR_add[5][9] ), .OUT(m1848) );
  XOR2 U3402 ( .A(\PR_mul[7][8] ), .B(\PR_add[5][8] ), .OUT(m1850) );
  XOR2 U3403 ( .A(m2322), .B(\PR_add[5][7] ), .OUT(m1852) );
  XOR2 U3404 ( .A(\PR_mul[7][6] ), .B(\PR_add[5][6] ), .OUT(m1854) );
  XOR2 U3405 ( .A(m2319), .B(\PR_add[5][5] ), .OUT(m1856) );
  XOR2 U3406 ( .A(\PR_mul[7][4] ), .B(\PR_add[5][4] ), .OUT(m1858) );
  XOR2 U3407 ( .A(m2316), .B(\PR_add[5][3] ), .OUT(m1860) );
  XOR2 U3408 ( .A(\PR_mul[7][2] ), .B(\PR_add[5][2] ), .OUT(m1862) );
  XOR2 U3409 ( .A(m2049), .B(\PR_add[5][1] ), .OUT(m2148) );
  XOR2 U3410 ( .A(m2056), .B(\PR_add[4][10] ), .OUT(m1864) );
  XOR2 U3411 ( .A(\PR_mul[6][9] ), .B(\PR_add[4][9] ), .OUT(m1866) );
  XOR2 U3412 ( .A(m2333), .B(\PR_add[4][8] ), .OUT(m1868) );
  XOR2 U3413 ( .A(\PR_mul[6][7] ), .B(\PR_add[4][7] ), .OUT(m1870) );
  XOR2 U3414 ( .A(m2330), .B(\PR_add[4][6] ), .OUT(m1872) );
  XOR2 U3415 ( .A(\PR_mul[6][5] ), .B(\PR_add[4][5] ), .OUT(m1874) );
  XOR2 U3416 ( .A(m2055), .B(\PR_add[4][4] ), .OUT(m2153) );
  XOR2 U3417 ( .A(m2062), .B(\PR_add[3][10] ), .OUT(m1876) );
  XOR2 U3418 ( .A(\PR_mul[5][9] ), .B(\PR_add[3][9] ), .OUT(m1878) );
  XOR2 U3419 ( .A(\PR_mul[5][8] ), .B(\PR_add[3][8] ), .OUT(m1880) );
  XOR2 U3420 ( .A(m2344), .B(\PR_add[3][7] ), .OUT(m1882) );
  XOR2 U3421 ( .A(\PR_mul[5][6] ), .B(\PR_add[3][6] ), .OUT(m1884) );
  XOR2 U3422 ( .A(m2341), .B(\PR_add[3][5] ), .OUT(m1886) );
  XOR2 U3423 ( .A(\PR_mul[5][4] ), .B(\PR_add[3][4] ), .OUT(m1888) );
  XOR2 U3424 ( .A(m2338), .B(\PR_add[3][3] ), .OUT(m1890) );
  XOR2 U3425 ( .A(\PR_mul[5][2] ), .B(\PR_add[3][2] ), .OUT(m1892) );
  XOR2 U3426 ( .A(m2061), .B(\PR_add[3][1] ), .OUT(m2158) );
  XOR2 U3427 ( .A(m2068), .B(\PR_add[2][9] ), .OUT(m1894) );
  XOR2 U3428 ( .A(\PR_mul[4][8] ), .B(\PR_add[2][8] ), .OUT(m1896) );
  XOR2 U3429 ( .A(m2354), .B(\PR_add[2][7] ), .OUT(m1898) );
  XOR2 U3430 ( .A(\PR_mul[4][6] ), .B(\PR_add[2][6] ), .OUT(m1900) );
  XOR2 U3431 ( .A(m2351), .B(\PR_add[2][5] ), .OUT(m1902) );
  XOR2 U3432 ( .A(\PR_mul[4][4] ), .B(\PR_add[2][4] ), .OUT(m1904) );
  XOR2 U3433 ( .A(m2067), .B(\PR_add[2][3] ), .OUT(m2163) );
  XOR2 U3434 ( .A(m2073), .B(\PR_add[1][11] ), .OUT(m1906) );
  XOR2 U3435 ( .A(\PR_mul[3][10] ), .B(\PR_add[1][10] ), .OUT(m1908) );
  XOR2 U3436 ( .A(m2366), .B(\PR_add[1][9] ), .OUT(m1910) );
  XOR2 U3437 ( .A(\PR_mul[3][8] ), .B(\PR_add[1][8] ), .OUT(m1912) );
  XOR2 U3438 ( .A(m2363), .B(\PR_add[1][7] ), .OUT(m1914) );
  XOR2 U3439 ( .A(\PR_mul[3][6] ), .B(\PR_add[1][6] ), .OUT(m1916) );
  XOR2 U3440 ( .A(m2360), .B(\PR_add[1][5] ), .OUT(m1918) );
  XOR2 U3441 ( .A(\PR_mul[3][4] ), .B(\PR_add[1][4] ), .OUT(m1920) );
  XOR2 U3442 ( .A(m2357), .B(\PR_add[1][3] ), .OUT(m1922) );
  XOR2 U3443 ( .A(\PR_mul[3][2] ), .B(\PR_add[1][2] ), .OUT(N150) );
  XOR2 U3444 ( .A(m2079), .B(\PR_add[0][11] ), .OUT(m1924) );
  XOR2 U3445 ( .A(\PR_mul[2][10] ), .B(\PR_add[0][10] ), .OUT(m1926) );
  XOR2 U3446 ( .A(m2380), .B(\PR_add[0][9] ), .OUT(m1928) );
  XOR2 U3447 ( .A(\PR_mul[2][8] ), .B(\PR_add[0][8] ), .OUT(m1930) );
  XOR2 U3448 ( .A(m2377), .B(\PR_add[0][7] ), .OUT(m1932) );
  XOR2 U3449 ( .A(\PR_mul[2][6] ), .B(\PR_add[0][6] ), .OUT(m1934) );
  XOR2 U3450 ( .A(m2374), .B(\PR_add[0][5] ), .OUT(m1936) );
  XOR2 U3451 ( .A(\PR_mul[2][4] ), .B(\PR_add[0][4] ), .OUT(m1938) );
  XOR2 U3452 ( .A(m2371), .B(\PR_add[0][3] ), .OUT(m1940) );
  XOR2 U3453 ( .A(\PR_mul[2][2] ), .B(\PR_add[0][2] ), .OUT(m1942) );
  XOR2 U3454 ( .A(m2078), .B(\PR_add[0][1] ), .OUT(m2170) );
  XOR2 U3455 ( .A(m1340), .B(\PR_mul[0][10] ), .OUT(m1944) );
  XOR2 U3456 ( .A(\PR_mul[1][9] ), .B(\PR_mul[0][9] ), .OUT(m1945) );
  XOR2 U3457 ( .A(m2388), .B(\PR_mul[0][8] ), .OUT(m1947) );
  XOR2 U3458 ( .A(\PR_mul[1][7] ), .B(\PR_mul[0][7] ), .OUT(m1949) );
  XOR2 U3459 ( .A(m2385), .B(\PR_mul[0][6] ), .OUT(m1951) );
  XOR2 U3460 ( .A(\PR_mul[1][5] ), .B(\PR_mul[0][5] ), .OUT(m1953) );
  XOR2 U3461 ( .A(m2081), .B(\PR_mul[0][4] ), .OUT(m2172) );
  INV U3462 ( .IN(m1345), .OUT(m2174) );
  INV U3463 ( .IN(m1347), .OUT(m2177) );
  INV U3464 ( .IN(m1349), .OUT(m2180) );
  INV U3465 ( .IN(m1956), .OUT(m1351) );
  INV U3466 ( .IN(m1354), .OUT(m1958) );
  INV U3467 ( .IN(m1357), .OUT(m1959) );
  INV U3468 ( .IN(m1360), .OUT(m2181) );
  INV U3469 ( .IN(m1362), .OUT(m2184) );
  INV U3470 ( .IN(m1369), .OUT(m1963) );
  INV U3471 ( .IN(m1372), .OUT(m1966) );
  INV U3472 ( .IN(m1378), .OUT(m2194) );
  INV U3473 ( .IN(m1381), .OUT(m2196) );
  INV U3474 ( .IN(m1383), .OUT(m2199) );
  INV U3475 ( .IN(m1385), .OUT(m2202) );
  INV U3476 ( .IN(m1974), .OUT(m1387) );
  INV U3477 ( .IN(m1390), .OUT(m1976) );
  INV U3478 ( .IN(m1393), .OUT(m1977) );
  INV U3479 ( .IN(m1396), .OUT(m2203) );
  INV U3480 ( .IN(m1398), .OUT(m2206) );
  INV U3481 ( .IN(m1405), .OUT(m1981) );
  INV U3482 ( .IN(m1408), .OUT(m1984) );
  INV U3483 ( .IN(m1414), .OUT(m2216) );
  INV U3484 ( .IN(m1417), .OUT(m2218) );
  INV U3485 ( .IN(m1419), .OUT(m2221) );
  INV U3486 ( .IN(m1421), .OUT(m2224) );
  INV U3487 ( .IN(m1992), .OUT(m1423) );
  INV U3488 ( .IN(m1426), .OUT(m1994) );
  INV U3489 ( .IN(m1429), .OUT(m1995) );
  INV U3490 ( .IN(m1432), .OUT(m2225) );
  INV U3491 ( .IN(m1434), .OUT(m2228) );
  INV U3492 ( .IN(m1441), .OUT(m1999) );
  INV U3493 ( .IN(m1444), .OUT(m2002) );
  INV U3494 ( .IN(m1450), .OUT(m2238) );
  INV U3495 ( .IN(m1453), .OUT(m2240) );
  INV U3496 ( .IN(m1455), .OUT(m2243) );
  INV U3497 ( .IN(m1457), .OUT(m2246) );
  INV U3498 ( .IN(\PR_add[12][13] ), .OUT(m2012) );
  INV U3499 ( .IN(m1472), .OUT(m2249) );
  INV U3500 ( .IN(m1474), .OUT(m2252) );
  INV U3501 ( .IN(m1476), .OUT(m2255) );
  INV U3502 ( .IN(m1478), .OUT(m2258) );
  INV U3503 ( .IN(m1488), .OUT(m2260) );
  INV U3504 ( .IN(m1490), .OUT(m2263) );
  INV U3505 ( .IN(m1492), .OUT(m2266) );
  INV U3506 ( .IN(m1494), .OUT(m2269) );
  INV U3507 ( .IN(m1496), .OUT(m2272) );
  INV U3508 ( .IN(m1506), .OUT(m2274) );
  INV U3509 ( .IN(m1508), .OUT(m2277) );
  INV U3510 ( .IN(m1510), .OUT(m2280) );
  INV U3511 ( .IN(\PR_add[9][14] ), .OUT(m2029) );
  INV U3512 ( .IN(m1522), .OUT(m2282) );
  INV U3513 ( .IN(m1524), .OUT(m2285) );
  INV U3514 ( .IN(m1526), .OUT(m2288) );
  INV U3515 ( .IN(m1528), .OUT(m2292) );
  INV U3516 ( .IN(m2291), .OUT(m1799) );
  INV U3517 ( .IN(m1529), .OUT(m2293) );
  INV U3518 ( .IN(\PR_add[8][14] ), .OUT(m2035) );
  INV U3519 ( .IN(m1541), .OUT(m2295) );
  INV U3520 ( .IN(m1543), .OUT(m2298) );
  INV U3521 ( .IN(m1545), .OUT(m2301) );
  INV U3522 ( .IN(\PR_add[7][13] ), .OUT(m2041) );
  INV U3523 ( .IN(m1560), .OUT(m2304) );
  INV U3524 ( .IN(m1562), .OUT(m2307) );
  INV U3525 ( .IN(m1564), .OUT(m2310) );
  INV U3526 ( .IN(m1566), .OUT(m2313) );
  INV U3527 ( .IN(m1576), .OUT(m2315) );
  INV U3528 ( .IN(m1578), .OUT(m2318) );
  INV U3529 ( .IN(m1580), .OUT(m2321) );
  INV U3530 ( .IN(m1582), .OUT(m2324) );
  INV U3531 ( .IN(m1584), .OUT(m2327) );
  INV U3532 ( .IN(m1594), .OUT(m2329) );
  INV U3533 ( .IN(m1596), .OUT(m2332) );
  INV U3534 ( .IN(m1598), .OUT(m2335) );
  INV U3535 ( .IN(\PR_add[4][14] ), .OUT(m2058) );
  INV U3536 ( .IN(m1610), .OUT(m2337) );
  INV U3537 ( .IN(m1612), .OUT(m2340) );
  INV U3538 ( .IN(m1614), .OUT(m2343) );
  INV U3539 ( .IN(m1616), .OUT(m2347) );
  INV U3540 ( .IN(m2346), .OUT(m1879) );
  INV U3541 ( .IN(m1617), .OUT(m2348) );
  INV U3542 ( .IN(\PR_add[3][14] ), .OUT(m2064) );
  INV U3543 ( .IN(m1629), .OUT(m2350) );
  INV U3544 ( .IN(m1631), .OUT(m2353) );
  INV U3545 ( .IN(m1633), .OUT(m2356) );
  INV U3546 ( .IN(\PR_add[2][13] ), .OUT(m2070) );
  INV U3547 ( .IN(m1648), .OUT(m2359) );
  INV U3548 ( .IN(m1650), .OUT(m2362) );
  INV U3549 ( .IN(m1652), .OUT(m2365) );
  INV U3550 ( .IN(m1654), .OUT(m2368) );
  INV U3551 ( .IN(m1664), .OUT(m2370) );
  INV U3552 ( .IN(m1666), .OUT(m2373) );
  INV U3553 ( .IN(m1668), .OUT(m2376) );
  INV U3554 ( .IN(m1670), .OUT(m2379) );
  INV U3555 ( .IN(m1672), .OUT(m2382) );
  INV U3556 ( .IN(m1675), .OUT(m2384) );
  INV U3557 ( .IN(m1677), .OUT(m2387) );
  INV U3558 ( .IN(m1679), .OUT(m2390) );
  INV U3559 ( .IN(\mult_83/ab[1][3] ), .OUT(m2082) );
  INV U3560 ( .IN(\mult_83/ab[2][2] ), .OUT(m2173) );
  INV U3561 ( .IN(\mult_83/ab[3][3] ), .OUT(m2175) );
  INV U3562 ( .IN(\mult_83/ab[4][2] ), .OUT(m2176) );
  INV U3563 ( .IN(\mult_83/ab[5][3] ), .OUT(m2178) );
  INV U3564 ( .IN(\mult_83/ab[6][2] ), .OUT(m2179) );
  INV U3565 ( .IN(\mult_80/ab[3][2] ), .OUT(m2186) );
  INV U3566 ( .IN(\mult_80/ab[4][1] ), .OUT(m2187) );
  INV U3567 ( .IN(\mult_80/ab[5][2] ), .OUT(m2191) );
  INV U3568 ( .IN(\mult_80/ab[6][1] ), .OUT(m2192) );
  INV U3569 ( .IN(\mult_77/ab[1][3] ), .OUT(m2091) );
  INV U3570 ( .IN(\mult_77/ab[2][2] ), .OUT(m2195) );
  INV U3571 ( .IN(\mult_77/ab[3][3] ), .OUT(m2197) );
  INV U3572 ( .IN(\mult_77/ab[4][2] ), .OUT(m2198) );
  INV U3573 ( .IN(\mult_77/ab[5][3] ), .OUT(m2200) );
  INV U3574 ( .IN(\mult_77/ab[6][2] ), .OUT(m2201) );
  INV U3575 ( .IN(\mult_74/ab[3][2] ), .OUT(m2208) );
  INV U3576 ( .IN(\mult_74/ab[4][1] ), .OUT(m2209) );
  INV U3577 ( .IN(\mult_74/ab[5][2] ), .OUT(m2213) );
  INV U3578 ( .IN(\mult_74/ab[6][1] ), .OUT(m2214) );
  INV U3579 ( .IN(\mult_72/ab[1][3] ), .OUT(m2100) );
  INV U3580 ( .IN(\mult_72/ab[2][2] ), .OUT(m2217) );
  INV U3581 ( .IN(\mult_72/ab[3][3] ), .OUT(m2219) );
  INV U3582 ( .IN(\mult_72/ab[4][2] ), .OUT(m2220) );
  INV U3583 ( .IN(\mult_72/ab[5][3] ), .OUT(m2222) );
  INV U3584 ( .IN(\mult_72/ab[6][2] ), .OUT(m2223) );
  INV U3585 ( .IN(\mult_69/ab[3][2] ), .OUT(m2230) );
  INV U3586 ( .IN(\mult_69/ab[4][1] ), .OUT(m2231) );
  INV U3587 ( .IN(\mult_69/ab[5][2] ), .OUT(m2235) );
  INV U3588 ( .IN(\mult_69/ab[6][1] ), .OUT(m2236) );
  INV U3589 ( .IN(\PR_mul[14][3] ), .OUT(m2112) );
  INV U3590 ( .IN(\PR_add[12][3] ), .OUT(m2239) );
  INV U3591 ( .IN(\PR_mul[14][5] ), .OUT(m2241) );
  INV U3592 ( .IN(\PR_add[12][5] ), .OUT(m2242) );
  INV U3593 ( .IN(\PR_mul[14][7] ), .OUT(m2244) );
  INV U3594 ( .IN(\PR_add[12][7] ), .OUT(m2245) );
  INV U3595 ( .IN(\PR_mul[13][3] ), .OUT(m2247) );
  INV U3596 ( .IN(\PR_add[11][3] ), .OUT(m2248) );
  INV U3597 ( .IN(\PR_mul[13][5] ), .OUT(m2250) );
  INV U3598 ( .IN(\PR_add[11][5] ), .OUT(m2251) );
  INV U3599 ( .IN(\PR_mul[13][7] ), .OUT(m2253) );
  INV U3600 ( .IN(\PR_add[11][7] ), .OUT(m2254) );
  INV U3601 ( .IN(\PR_mul[13][9] ), .OUT(m2256) );
  INV U3602 ( .IN(\PR_add[11][9] ), .OUT(m2257) );
  INV U3603 ( .IN(\PR_mul[12][1] ), .OUT(m2122) );
  INV U3604 ( .IN(\PR_add[10][1] ), .OUT(m2259) );
  INV U3605 ( .IN(\PR_mul[12][3] ), .OUT(m2261) );
  INV U3606 ( .IN(\PR_add[10][3] ), .OUT(m2262) );
  INV U3607 ( .IN(\PR_mul[12][5] ), .OUT(m2264) );
  INV U3608 ( .IN(\PR_add[10][5] ), .OUT(m2265) );
  INV U3609 ( .IN(\PR_mul[12][7] ), .OUT(m2267) );
  INV U3610 ( .IN(\PR_add[10][7] ), .OUT(m2268) );
  INV U3611 ( .IN(\PR_mul[12][9] ), .OUT(m2270) );
  INV U3612 ( .IN(\PR_add[10][9] ), .OUT(m2271) );
  INV U3613 ( .IN(\PR_mul[11][4] ), .OUT(m2127) );
  INV U3614 ( .IN(\PR_add[9][4] ), .OUT(m2273) );
  INV U3615 ( .IN(\PR_mul[11][6] ), .OUT(m2275) );
  INV U3616 ( .IN(\PR_add[9][6] ), .OUT(m2276) );
  INV U3617 ( .IN(\PR_mul[11][8] ), .OUT(m2278) );
  INV U3618 ( .IN(\PR_add[9][8] ), .OUT(m2279) );
  INV U3619 ( .IN(\PR_mul[10][1] ), .OUT(m2132) );
  INV U3620 ( .IN(\PR_add[8][1] ), .OUT(m2281) );
  INV U3621 ( .IN(\PR_mul[10][3] ), .OUT(m2283) );
  INV U3622 ( .IN(\PR_add[8][3] ), .OUT(m2284) );
  INV U3623 ( .IN(\PR_mul[10][5] ), .OUT(m2286) );
  INV U3624 ( .IN(\PR_add[8][5] ), .OUT(m2287) );
  INV U3625 ( .IN(\PR_mul[10][7] ), .OUT(m2289) );
  INV U3626 ( .IN(\PR_add[8][7] ), .OUT(m2290) );
  INV U3627 ( .IN(\PR_mul[9][3] ), .OUT(m2137) );
  INV U3628 ( .IN(\PR_add[7][3] ), .OUT(m2294) );
  INV U3629 ( .IN(\PR_mul[9][5] ), .OUT(m2296) );
  INV U3630 ( .IN(\PR_add[7][5] ), .OUT(m2297) );
  INV U3631 ( .IN(\PR_mul[9][7] ), .OUT(m2299) );
  INV U3632 ( .IN(\PR_add[7][7] ), .OUT(m2300) );
  INV U3633 ( .IN(\PR_mul[8][3] ), .OUT(m2302) );
  INV U3634 ( .IN(\PR_add[6][3] ), .OUT(m2303) );
  INV U3635 ( .IN(\PR_mul[8][5] ), .OUT(m2305) );
  INV U3636 ( .IN(\PR_add[6][5] ), .OUT(m2306) );
  INV U3637 ( .IN(\PR_mul[8][7] ), .OUT(m2308) );
  INV U3638 ( .IN(\PR_add[6][7] ), .OUT(m2309) );
  INV U3639 ( .IN(\PR_mul[8][9] ), .OUT(m2311) );
  INV U3640 ( .IN(\PR_add[6][9] ), .OUT(m2312) );
  INV U3641 ( .IN(\PR_mul[7][1] ), .OUT(m2147) );
  INV U3642 ( .IN(\PR_add[5][1] ), .OUT(m2314) );
  INV U3643 ( .IN(\PR_mul[7][3] ), .OUT(m2316) );
  INV U3644 ( .IN(\PR_add[5][3] ), .OUT(m2317) );
  INV U3645 ( .IN(\PR_mul[7][5] ), .OUT(m2319) );
  INV U3646 ( .IN(\PR_add[5][5] ), .OUT(m2320) );
  INV U3647 ( .IN(\PR_mul[7][7] ), .OUT(m2322) );
  INV U3648 ( .IN(\PR_add[5][7] ), .OUT(m2323) );
  INV U3649 ( .IN(\PR_mul[7][9] ), .OUT(m2325) );
  INV U3650 ( .IN(\PR_add[5][9] ), .OUT(m2326) );
  INV U3651 ( .IN(\PR_mul[6][4] ), .OUT(m2152) );
  INV U3652 ( .IN(\PR_add[4][4] ), .OUT(m2328) );
  INV U3653 ( .IN(\PR_mul[6][6] ), .OUT(m2330) );
  INV U3654 ( .IN(\PR_add[4][6] ), .OUT(m2331) );
  INV U3655 ( .IN(\PR_mul[6][8] ), .OUT(m2333) );
  INV U3656 ( .IN(\PR_add[4][8] ), .OUT(m2334) );
  INV U3657 ( .IN(\PR_mul[5][1] ), .OUT(m2157) );
  INV U3658 ( .IN(\PR_add[3][1] ), .OUT(m2336) );
  INV U3659 ( .IN(\PR_mul[5][3] ), .OUT(m2338) );
  INV U3660 ( .IN(\PR_add[3][3] ), .OUT(m2339) );
  INV U3661 ( .IN(\PR_mul[5][5] ), .OUT(m2341) );
  INV U3662 ( .IN(\PR_add[3][5] ), .OUT(m2342) );
  INV U3663 ( .IN(\PR_mul[5][7] ), .OUT(m2344) );
  INV U3664 ( .IN(\PR_add[3][7] ), .OUT(m2345) );
  INV U3665 ( .IN(\PR_mul[4][3] ), .OUT(m2162) );
  INV U3666 ( .IN(\PR_add[2][3] ), .OUT(m2349) );
  INV U3667 ( .IN(\PR_mul[4][5] ), .OUT(m2351) );
  INV U3668 ( .IN(\PR_add[2][5] ), .OUT(m2352) );
  INV U3669 ( .IN(\PR_mul[4][7] ), .OUT(m2354) );
  INV U3670 ( .IN(\PR_add[2][7] ), .OUT(m2355) );
  INV U3671 ( .IN(\PR_mul[3][3] ), .OUT(m2357) );
  INV U3672 ( .IN(\PR_add[1][3] ), .OUT(m2358) );
  INV U3673 ( .IN(\PR_mul[3][5] ), .OUT(m2360) );
  INV U3674 ( .IN(\PR_add[1][5] ), .OUT(m2361) );
  INV U3675 ( .IN(\PR_mul[3][7] ), .OUT(m2363) );
  INV U3676 ( .IN(\PR_add[1][7] ), .OUT(m2364) );
  INV U3677 ( .IN(\PR_mul[3][9] ), .OUT(m2366) );
  INV U3678 ( .IN(\PR_add[1][9] ), .OUT(m2367) );
  INV U3679 ( .IN(\PR_mul[2][1] ), .OUT(m2169) );
  INV U3680 ( .IN(\PR_add[0][1] ), .OUT(m2369) );
  INV U3681 ( .IN(\PR_mul[2][3] ), .OUT(m2371) );
  INV U3682 ( .IN(\PR_add[0][3] ), .OUT(m2372) );
  INV U3683 ( .IN(\PR_mul[2][5] ), .OUT(m2374) );
  INV U3684 ( .IN(\PR_add[0][5] ), .OUT(m2375) );
  INV U3685 ( .IN(\PR_mul[2][7] ), .OUT(m2377) );
  INV U3686 ( .IN(\PR_add[0][7] ), .OUT(m2378) );
  INV U3687 ( .IN(\PR_mul[2][9] ), .OUT(m2380) );
  INV U3688 ( .IN(\PR_add[0][9] ), .OUT(m2381) );
  INV U3689 ( .IN(\PR_mul[1][4] ), .OUT(m2171) );
  INV U3690 ( .IN(\PR_mul[0][4] ), .OUT(m2383) );
  INV U3691 ( .IN(\PR_mul[1][6] ), .OUT(m2385) );
  INV U3692 ( .IN(\PR_mul[0][6] ), .OUT(m2386) );
  INV U3693 ( .IN(\PR_mul[1][8] ), .OUT(m2388) );
  INV U3694 ( .IN(\PR_mul[0][8] ), .OUT(m2389) );
  INV U3695 ( .IN(m1962), .OUT(m1371) );
  INV U3696 ( .IN(m1965), .OUT(m1375) );
  INV U3697 ( .IN(m1980), .OUT(m1407) );
  INV U3698 ( .IN(m1983), .OUT(m1411) );
  INV U3699 ( .IN(m1998), .OUT(m1443) );
  INV U3700 ( .IN(m2001), .OUT(m1447) );
  INV U3701 ( .IN(m1350), .OUT(m1957) );
  INV U3702 ( .IN(m1364), .OUT(m2189) );
  INV U3703 ( .IN(m1366), .OUT(m2193) );
  INV U3704 ( .IN(\mult_80/ab[2][0] ), .OUT(m1368) );
  INV U3705 ( .IN(m2393), .OUT(m1972) );
  INV U3706 ( .IN(m2396), .OUT(m1337) );
  INV U3707 ( .IN(m1386), .OUT(m1975) );
  INV U3708 ( .IN(m1400), .OUT(m2211) );
  INV U3709 ( .IN(m1402), .OUT(m2215) );
  INV U3710 ( .IN(\mult_74/ab[2][0] ), .OUT(m1404) );
  INV U3711 ( .IN(m2400), .OUT(m1990) );
  INV U3712 ( .IN(m2403), .OUT(m1329) );
  INV U3713 ( .IN(m1422), .OUT(m1993) );
  INV U3714 ( .IN(m1436), .OUT(m2233) );
  INV U3715 ( .IN(m1438), .OUT(m2237) );
  INV U3716 ( .IN(\mult_69/ab[2][0] ), .OUT(m1440) );
  INV U3717 ( .IN(m2407), .OUT(m2008) );
  INV U3718 ( .IN(m2410), .OUT(m1321) );
  INV U3719 ( .IN(m2109), .OUT(N385) );
  INV U3720 ( .IN(m2110), .OUT(N383) );
  INV U3721 ( .IN(m2111), .OUT(N379) );
  INV U3722 ( .IN(m2114), .OUT(N365) );
  INV U3723 ( .IN(m2116), .OUT(N361) );
  INV U3724 ( .IN(m2119), .OUT(N345) );
  INV U3725 ( .IN(m2121), .OUT(N341) );
  INV U3726 ( .IN(m2124), .OUT(N327) );
  INV U3727 ( .IN(m2125), .OUT(N324) );
  INV U3728 ( .IN(m2126), .OUT(N320) );
  INV U3729 ( .IN(m2129), .OUT(N307) );
  INV U3730 ( .IN(m2130), .OUT(N304) );
  INV U3731 ( .IN(m2131), .OUT(N300) );
  INV U3732 ( .IN(m2134), .OUT(N285) );
  INV U3733 ( .IN(m2135), .OUT(N283) );
  INV U3734 ( .IN(m2136), .OUT(N279) );
  INV U3735 ( .IN(m2139), .OUT(N265) );
  INV U3736 ( .IN(m2141), .OUT(N261) );
  INV U3737 ( .IN(m2144), .OUT(N245) );
  INV U3738 ( .IN(m2146), .OUT(N241) );
  INV U3739 ( .IN(m2149), .OUT(N227) );
  INV U3740 ( .IN(m2150), .OUT(N224) );
  INV U3741 ( .IN(m2151), .OUT(N220) );
  INV U3742 ( .IN(m2154), .OUT(N207) );
  INV U3743 ( .IN(m2155), .OUT(N204) );
  INV U3744 ( .IN(m2156), .OUT(N200) );
  INV U3745 ( .IN(m2159), .OUT(N185) );
  INV U3746 ( .IN(m2160), .OUT(N183) );
  INV U3747 ( .IN(m2161), .OUT(N179) );
  INV U3748 ( .IN(m2164), .OUT(N165) );
  INV U3749 ( .IN(m2166), .OUT(N161) );
  INV U3750 ( .IN(\mult_82/A1[0] ), .OUT(m2412) );
  INV U3751 ( .IN(m2413), .OUT(N86) );
  INV U3752 ( .IN(\mult_82/A1[1] ), .OUT(m2414) );
  INV U3753 ( .IN(m2415), .OUT(N87) );
  INV U3754 ( .IN(\mult_82/A1[2] ), .OUT(m2416) );
  INV U3755 ( .IN(m2417), .OUT(N88) );
  INV U3756 ( .IN(\mult_82/A1[3] ), .OUT(m2418) );
  INV U3757 ( .IN(m2419), .OUT(N89) );
  INV U3758 ( .IN(\mult_82/A1[4] ), .OUT(m2420) );
  INV U3759 ( .IN(m2421), .OUT(N90) );
  INV U3760 ( .IN(\mult_82/A1[5] ), .OUT(m2422) );
  INV U3761 ( .IN(m2423), .OUT(N91) );
  INV U3762 ( .IN(\mult_82/A1[6] ), .OUT(m2424) );
  INV U3763 ( .IN(m2425), .OUT(N92) );
  INV U3764 ( .IN(\mult_82/A1[7] ), .OUT(m2426) );
  INV U3765 ( .IN(\mult_82/A2[7] ), .OUT(m2427) );
  INV U3766 ( .IN(\mult_82/FS_1/G_n_int[0][1][3] ), .OUT(
        \mult_82/FS_1/G[0][1][3] ) );
  INV U3767 ( .IN(m2428), .OUT(N93) );
  INV U3768 ( .IN(m2429), .OUT(\mult_82/FS_1/G[1][0][1] ) );
  INV U3769 ( .IN(\mult_82/A1[8] ), .OUT(m2430) );
  INV U3770 ( .IN(m2431), .OUT(\mult_82/FS_1/PG_int[0][2][0] ) );
  INV U3771 ( .IN(m2432), .OUT(N95) );
  INV U3772 ( .IN(m2433), .OUT(\mult_82/FS_1/C[1][2][0] ) );
  INV U3773 ( .IN(\mult_69/A1[0] ), .OUT(m2434) );
  INV U3774 ( .IN(m2435), .OUT(N5) );
  INV U3775 ( .IN(\mult_69/A1[1] ), .OUT(m2436) );
  INV U3776 ( .IN(m2437), .OUT(N6) );
  INV U3777 ( .IN(\mult_69/A1[2] ), .OUT(m2438) );
  INV U3778 ( .IN(m2439), .OUT(N7) );
  INV U3779 ( .IN(\mult_69/A1[3] ), .OUT(m2440) );
  INV U3780 ( .IN(m2441), .OUT(N8) );
  INV U3781 ( .IN(\mult_69/A1[4] ), .OUT(m2442) );
  INV U3782 ( .IN(m2443), .OUT(N9) );
  INV U3783 ( .IN(\mult_69/A1[5] ), .OUT(m2444) );
  INV U3784 ( .IN(m2445), .OUT(N10) );
  INV U3785 ( .IN(\mult_69/A1[6] ), .OUT(m2446) );
  INV U3786 ( .IN(m2447), .OUT(N11) );
  INV U3787 ( .IN(\mult_69/A1[7] ), .OUT(m2448) );
  INV U3788 ( .IN(\mult_69/A2[7] ), .OUT(m2449) );
  INV U3789 ( .IN(\mult_69/FS_1/G_n_int[0][1][3] ), .OUT(
        \mult_69/FS_1/G[0][1][3] ) );
  INV U3790 ( .IN(m2450), .OUT(N12) );
  INV U3791 ( .IN(m2451), .OUT(\mult_69/FS_1/G[1][0][1] ) );
  INV U3792 ( .IN(\mult_69/A2[8] ), .OUT(m2452) );
  INV U3793 ( .IN(m2453), .OUT(\mult_69/FS_1/PG_int[0][2][0] ) );
  INV U3794 ( .IN(m2454), .OUT(\mult_69/FS_1/C[1][2][0] ) );
  INV U3795 ( .IN(\mult_71/A1[0] ), .OUT(m2455) );
  INV U3796 ( .IN(m2456), .OUT(N16) );
  INV U3797 ( .IN(\mult_71/A1[1] ), .OUT(m2457) );
  INV U3798 ( .IN(m2458), .OUT(N17) );
  INV U3799 ( .IN(\mult_71/A1[2] ), .OUT(m2459) );
  INV U3800 ( .IN(m2460), .OUT(N18) );
  INV U3801 ( .IN(\mult_71/A1[3] ), .OUT(m2461) );
  INV U3802 ( .IN(m2462), .OUT(N19) );
  INV U3803 ( .IN(\mult_71/A1[4] ), .OUT(m2463) );
  INV U3804 ( .IN(m2464), .OUT(N20) );
  INV U3805 ( .IN(\mult_71/A1[5] ), .OUT(m2465) );
  INV U3806 ( .IN(m2466), .OUT(N21) );
  INV U3807 ( .IN(\mult_71/A1[6] ), .OUT(m2467) );
  INV U3808 ( .IN(m2468), .OUT(N22) );
  INV U3809 ( .IN(\mult_71/A1[7] ), .OUT(m2469) );
  INV U3810 ( .IN(\mult_71/A2[7] ), .OUT(m2470) );
  INV U3811 ( .IN(\mult_71/FS_1/G_n_int[0][1][3] ), .OUT(
        \mult_71/FS_1/G[0][1][3] ) );
  INV U3812 ( .IN(m2471), .OUT(N23) );
  INV U3813 ( .IN(m2472), .OUT(\mult_71/FS_1/G[1][0][1] ) );
  INV U3814 ( .IN(\mult_71/A1[8] ), .OUT(m2473) );
  INV U3815 ( .IN(m2474), .OUT(\mult_71/FS_1/PG_int[0][2][0] ) );
  INV U3816 ( .IN(m2475), .OUT(N25) );
  INV U3817 ( .IN(m2476), .OUT(\mult_71/FS_1/C[1][2][0] ) );
  INV U3818 ( .IN(\mult_72/A1[0] ), .OUT(m2477) );
  INV U3819 ( .IN(m2478), .OUT(N28) );
  INV U3820 ( .IN(\mult_72/A1[1] ), .OUT(m2479) );
  INV U3821 ( .IN(m2480), .OUT(N29) );
  INV U3822 ( .IN(\mult_72/A1[2] ), .OUT(m2481) );
  INV U3823 ( .IN(m2482), .OUT(N30) );
  INV U3824 ( .IN(\mult_72/A1[3] ), .OUT(m2483) );
  INV U3825 ( .IN(m2484), .OUT(N31) );
  INV U3826 ( .IN(\mult_72/A1[4] ), .OUT(m2485) );
  INV U3827 ( .IN(m2486), .OUT(N32) );
  INV U3828 ( .IN(\mult_72/A1[5] ), .OUT(m2487) );
  INV U3829 ( .IN(m2488), .OUT(N33) );
  INV U3830 ( .IN(\mult_72/A1[6] ), .OUT(m2489) );
  INV U3831 ( .IN(m2490), .OUT(N34) );
  INV U3832 ( .IN(\mult_72/A1[7] ), .OUT(m2491) );
  INV U3833 ( .IN(m2492), .OUT(N35) );
  INV U3834 ( .IN(\mult_72/A1[8] ), .OUT(m2493) );
  INV U3835 ( .IN(m2494), .OUT(N36) );
  INV U3836 ( .IN(\mult_72/A2[9] ), .OUT(m2495) );
  INV U3837 ( .IN(m2496), .OUT(N37) );
  INV U3838 ( .IN(\mult_74/A1[0] ), .OUT(m2497) );
  INV U3839 ( .IN(m2498), .OUT(N40) );
  INV U3840 ( .IN(\mult_74/A1[1] ), .OUT(m2499) );
  INV U3841 ( .IN(m2500), .OUT(N41) );
  INV U3842 ( .IN(\mult_74/A1[2] ), .OUT(m2501) );
  INV U3843 ( .IN(m2502), .OUT(N42) );
  INV U3844 ( .IN(\mult_74/A1[3] ), .OUT(m2503) );
  INV U3845 ( .IN(m2504), .OUT(N43) );
  INV U3846 ( .IN(\mult_74/A1[4] ), .OUT(m2505) );
  INV U3847 ( .IN(m2506), .OUT(N44) );
  INV U3848 ( .IN(\mult_74/A1[5] ), .OUT(m2507) );
  INV U3849 ( .IN(m2508), .OUT(N45) );
  INV U3850 ( .IN(\mult_74/A1[6] ), .OUT(m2509) );
  INV U3851 ( .IN(m2510), .OUT(N46) );
  INV U3852 ( .IN(\mult_74/A1[7] ), .OUT(m2511) );
  INV U3853 ( .IN(\mult_74/A2[7] ), .OUT(m2512) );
  INV U3854 ( .IN(\mult_74/FS_1/G_n_int[0][1][3] ), .OUT(
        \mult_74/FS_1/G[0][1][3] ) );
  INV U3855 ( .IN(m2513), .OUT(N47) );
  INV U3856 ( .IN(m2514), .OUT(\mult_74/FS_1/G[1][0][1] ) );
  INV U3857 ( .IN(\mult_74/A2[8] ), .OUT(m2515) );
  INV U3858 ( .IN(m2516), .OUT(\mult_74/FS_1/PG_int[0][2][0] ) );
  INV U3859 ( .IN(m2517), .OUT(\mult_74/FS_1/C[1][2][0] ) );
  INV U3860 ( .IN(\mult_76/A1[0] ), .OUT(m2518) );
  INV U3861 ( .IN(m2519), .OUT(N51) );
  INV U3862 ( .IN(\mult_76/A1[1] ), .OUT(m2520) );
  INV U3863 ( .IN(m2521), .OUT(N52) );
  INV U3864 ( .IN(\mult_76/A1[2] ), .OUT(m2522) );
  INV U3865 ( .IN(m2523), .OUT(N53) );
  INV U3866 ( .IN(\mult_76/A1[3] ), .OUT(m2524) );
  INV U3867 ( .IN(m2525), .OUT(N54) );
  INV U3868 ( .IN(\mult_76/A1[4] ), .OUT(m2526) );
  INV U3869 ( .IN(m2527), .OUT(N55) );
  INV U3870 ( .IN(\mult_76/A1[5] ), .OUT(m2528) );
  INV U3871 ( .IN(m2529), .OUT(N56) );
  INV U3872 ( .IN(\mult_76/A1[6] ), .OUT(m2530) );
  INV U3873 ( .IN(m2531), .OUT(N57) );
  INV U3874 ( .IN(\mult_76/A1[7] ), .OUT(m2532) );
  INV U3875 ( .IN(\mult_76/A2[7] ), .OUT(m2533) );
  INV U3876 ( .IN(\mult_76/FS_1/G_n_int[0][1][3] ), .OUT(
        \mult_76/FS_1/G[0][1][3] ) );
  INV U3877 ( .IN(m2534), .OUT(N58) );
  INV U3878 ( .IN(m2535), .OUT(\mult_76/FS_1/G[1][0][1] ) );
  INV U3879 ( .IN(\mult_76/A1[8] ), .OUT(m2536) );
  INV U3880 ( .IN(m2537), .OUT(\mult_76/FS_1/PG_int[0][2][0] ) );
  INV U3881 ( .IN(m2538), .OUT(N60) );
  INV U3882 ( .IN(m2539), .OUT(\mult_76/FS_1/C[1][2][0] ) );
  INV U3883 ( .IN(\mult_77/A1[0] ), .OUT(m2540) );
  INV U3884 ( .IN(m2541), .OUT(N63) );
  INV U3885 ( .IN(\mult_77/A1[1] ), .OUT(m2542) );
  INV U3886 ( .IN(m2543), .OUT(N64) );
  INV U3887 ( .IN(\mult_77/A1[2] ), .OUT(m2544) );
  INV U3888 ( .IN(m2545), .OUT(N65) );
  INV U3889 ( .IN(\mult_77/A1[3] ), .OUT(m2546) );
  INV U3890 ( .IN(m2547), .OUT(N66) );
  INV U3891 ( .IN(\mult_77/A1[4] ), .OUT(m2548) );
  INV U3892 ( .IN(m2549), .OUT(N67) );
  INV U3893 ( .IN(\mult_77/A1[5] ), .OUT(m2550) );
  INV U3894 ( .IN(m2551), .OUT(N68) );
  INV U3895 ( .IN(\mult_77/A1[6] ), .OUT(m2552) );
  INV U3896 ( .IN(m2553), .OUT(N69) );
  INV U3897 ( .IN(\mult_77/A1[7] ), .OUT(m2554) );
  INV U3898 ( .IN(m2555), .OUT(N70) );
  INV U3899 ( .IN(\mult_77/A1[8] ), .OUT(m2556) );
  INV U3900 ( .IN(m2557), .OUT(N71) );
  INV U3901 ( .IN(\mult_77/A2[9] ), .OUT(m2558) );
  INV U3902 ( .IN(m2559), .OUT(N72) );
  INV U3903 ( .IN(\mult_80/A1[0] ), .OUT(m2560) );
  INV U3904 ( .IN(m2561), .OUT(N75) );
  INV U3905 ( .IN(\mult_80/A1[1] ), .OUT(m2562) );
  INV U3906 ( .IN(m2563), .OUT(N76) );
  INV U3907 ( .IN(\mult_80/A1[2] ), .OUT(m2564) );
  INV U3908 ( .IN(m2565), .OUT(N77) );
  INV U3909 ( .IN(\mult_80/A1[3] ), .OUT(m2566) );
  INV U3910 ( .IN(m2567), .OUT(N78) );
  INV U3911 ( .IN(\mult_80/A1[4] ), .OUT(m2568) );
  INV U3912 ( .IN(m2569), .OUT(N79) );
  INV U3913 ( .IN(\mult_80/A1[5] ), .OUT(m2570) );
  INV U3914 ( .IN(m2571), .OUT(N80) );
  INV U3915 ( .IN(\mult_80/A1[6] ), .OUT(m2572) );
  INV U3916 ( .IN(m2573), .OUT(N81) );
  INV U3917 ( .IN(\mult_80/A1[7] ), .OUT(m2574) );
  INV U3918 ( .IN(\mult_80/A2[7] ), .OUT(m2575) );
  INV U3919 ( .IN(\mult_80/FS_1/G_n_int[0][1][3] ), .OUT(
        \mult_80/FS_1/G[0][1][3] ) );
  INV U3920 ( .IN(m2576), .OUT(N82) );
  INV U3921 ( .IN(m2577), .OUT(\mult_80/FS_1/G[1][0][1] ) );
  INV U3922 ( .IN(\mult_80/A2[8] ), .OUT(m2578) );
  INV U3923 ( .IN(m2579), .OUT(\mult_80/FS_1/PG_int[0][2][0] ) );
  INV U3924 ( .IN(m2580), .OUT(\mult_80/FS_1/C[1][2][0] ) );
  INV U3925 ( .IN(\mult_83/A1[0] ), .OUT(m2581) );
  INV U3926 ( .IN(m2582), .OUT(N98) );
  INV U3927 ( .IN(\mult_83/A1[1] ), .OUT(m2583) );
  INV U3928 ( .IN(m2584), .OUT(N99) );
  INV U3929 ( .IN(\mult_83/A1[2] ), .OUT(m2585) );
  INV U3930 ( .IN(m2586), .OUT(N100) );
  INV U3931 ( .IN(\mult_83/A1[3] ), .OUT(m2587) );
  INV U3932 ( .IN(m2588), .OUT(N101) );
  INV U3933 ( .IN(\mult_83/A1[4] ), .OUT(m2589) );
  INV U3934 ( .IN(m2590), .OUT(N102) );
  INV U3935 ( .IN(\mult_83/A1[5] ), .OUT(m2591) );
  INV U3936 ( .IN(m2592), .OUT(N103) );
  INV U3937 ( .IN(\mult_83/A1[6] ), .OUT(m2593) );
  INV U3938 ( .IN(m2594), .OUT(N104) );
  INV U3939 ( .IN(\mult_83/A1[7] ), .OUT(m2595) );
  INV U3940 ( .IN(m2596), .OUT(N105) );
  INV U3941 ( .IN(\mult_83/A1[8] ), .OUT(m2597) );
  INV U3942 ( .IN(m2598), .OUT(N106) );
  INV U3943 ( .IN(\mult_83/A2[9] ), .OUT(m2599) );
  INV U3944 ( .IN(m2600), .OUT(N107) );
endmodule

