* File: inv.pex.sp
* Created: Fri Oct 11 03:43:08 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.include "inv.pex.sp.pex"
.subckt inv  GND! OUT VDD! IN
* 
* IN	IN
* VDD!	VDD!
* OUT	OUT
* GND!	GND!
XD0_noxref N_GND!_D0_noxref_pos N_VDD!_D0_noxref_neg DIODENWX  AREA=2.9315e-12
+ PERIM=7.53e-06
XMMN0 N_OUT_MMN0_d N_IN_MMN0_g N_GND!_MMN0_s N_GND!_D0_noxref_pos NFET L=6.5e-08
+ W=1.7e-06 AD=4.913e-13 AS=4.182e-13 PD=3.978e-06 PS=3.892e-06 NRD=0.0970588
+ NRS=0.0888235 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=2.46e-07
+ SB=2.89e-07 SD=0 PANW1=0 PANW2=2.47e-15 PANW3=3.25e-15 PANW4=3.25e-15
+ PANW5=3.25e-15 PANW6=6.5e-15 PANW7=1.3e-14 PANW8=1.3e-14 PANW9=2.6e-14
+ PANW10=3.9e-14
XMMP0 N_OUT_MMP0_d N_IN_MMP0_g N_VDD!_MMP0_s N_VDD!_D0_noxref_neg PFET L=6.5e-08
+ W=1.8e-06 AD=5.004e-13 AS=4.626e-13 PD=4.156e-06 PS=4.114e-06 NRD=0.0919444
+ NRS=0.0926389 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=2.57e-07
+ SB=2.78e-07 SD=0 PANW1=0 PANW2=2.405e-15 PANW3=3.25e-15 PANW4=3.25e-15
+ PANW5=3.25e-15 PANW6=2.4362e-13 PANW7=2.6e-14 PANW8=2.6e-14 PANW9=5.2e-14
+ PANW10=7.8e-14
*
.include "inv.pex.sp.INV.pxi"
*
.ends
*
*
