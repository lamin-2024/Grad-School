* File: OAI12.pex.sp
* Created: Sat Nov  2 21:52:30 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.include "OAI12.pex.sp.pex"
.subckt OAI12  OUT VSS VDD VA VC VB
* 
* VB	VB
* VC	VC
* VA	VA
* VDD	VDD
* VSS	VSS
* OUT	OUT
XD0_noxref N_VSS_D0_noxref_pos N_VDD_D0_noxref_neg DIODENWX  AREA=9.48582e-12
+ PERIM=1.232e-05
XMMN0 N_OUT_MMN0_d N_VA_MMN0_g N_NET23_MMN0_s N_VSS_D0_noxref_pos NFET
+ L=6.2e-08 W=1.7e-06 AD=7.684e-13 AS=6.528e-13 PD=4.304e-06 PS=2.468e-06
+ NRD=0.133529 NRS=0.337059 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=4.52e-07 SB=1.793e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=6.2e-17
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=2.48e-14 PANW10=3.72e-14
XMMN4 N_NET23_MMN0_s N_VC_MMN4_g N_VSS_MMN4_s N_VSS_D0_noxref_pos NFET
+ L=6.2e-08 W=1.7e-06 AD=6.528e-13 AS=3.825e-13 PD=2.468e-06 PS=2.15e-06
+ NRD=0.114706 NRS=0.132353 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=1.282e-06 SB=9.63e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=6.2e-17
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=2.48e-14 PANW10=3.72e-14
XMMN1 N_NET23_MMN1_d N_VB_MMN1_g N_VSS_MMN4_s N_VSS_D0_noxref_pos NFET
+ L=6.2e-08 W=1.7e-06 AD=7.667e-13 AS=3.825e-13 PD=4.302e-06 PS=2.15e-06
+ NRD=0.132353 NRS=0.132353 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=1.794e-06 SB=4.51e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=6.2e-17
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=2.48e-14 PANW10=3.72e-14
XMMP0 N_OUT_MMP0_d N_VA_MMP0_g N_VDD_MMP0_s N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=1.8e-06 AD=6.912e-13 AS=8.136e-13 PD=2.568e-06 PS=4.504e-06 NRD=0.213333
+ NRS=0.126111 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=4.52e-07
+ SB=1.793e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=1.674e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.34478e-13 PANW9=4.96e-14 PANW10=7.44e-14
XMMP1 N_OUT_MMP0_d N_VC_MMP1_g NET8 N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=1.8e-06 AD=6.912e-13 AS=4.05e-13 PD=2.568e-06 PS=2.25e-06 NRD=0.213333
+ NRS=0.125 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.282e-06
+ SB=9.63e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=1.674e-15 PANW6=6.2e-15
+ PANW7=1.24e-14 PANW8=2.2878e-14 PANW9=1.612e-13 PANW10=1.86e-13
XMMP4 NET8 N_VB_MMP4_g N_VDD_MMP4_s N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=1.8e-06 AD=4.05e-13 AS=8.118e-13 PD=2.25e-06 PS=4.502e-06 NRD=0.125
+ NRS=0.125556 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.794e-06
+ SB=4.51e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=1.674e-15 PANW6=6.2e-15
+ PANW7=1.24e-14 PANW8=1.34478e-13 PANW9=4.96e-14 PANW10=7.44e-14
*
.include "OAI12.pex.sp.OAI12.pxi"
*
.ends
*
*
