* File: OAI12.pex.sp
* Created: Mon Dec  2 11:00:25 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.include "OAI12.pex.sp.pex"
.subckt OAI12  OUT VSS VDD A C B
* 
* B	B
* C	C
* A	A
* VDD	VDD
* VSS	VSS
* OUT	OUT
XD0_noxref N_VSS_D0_noxref_pos N_VDD_D0_noxref_neg DIODENWX  AREA=1.17925e-11
+ PERIM=1.3826e-05
XMMN0 N_OUT_MMN0_d N_A_MMN0_g N_NET23_MMN0_s N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=1.7e-06 AD=7.684e-13 AS=6.6215e-13 PD=4.304e-06 PS=2.479e-06 NRD=0.133529
+ NRS=0.339412 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=4.52e-07
+ SB=1.812e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=3.348e-15 PANW9=2.48e-14 PANW10=3.72e-14
XMMN4 N_NET23_MMN0_s N_C_MMN4_g N_VSS_MMN4_s N_VSS_D0_noxref_pos NFET
+ L=6.2e-08 W=1.7e-06 AD=6.6215e-13 AS=3.893e-13 PD=2.479e-06 PS=2.158e-06
+ NRD=0.118824 NRS=0.132353 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=1.293e-06 SB=9.71e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=0 PANW8=3.348e-15 PANW9=2.48e-14 PANW10=3.72e-14
XMMN1 N_NET23_MMN1_d N_B_MMN1_g N_VSS_MMN4_s N_VSS_D0_noxref_pos NFET
+ L=6.2e-08 W=1.7e-06 AD=7.667e-13 AS=3.893e-13 PD=4.302e-06 PS=2.158e-06
+ NRD=0.132353 NRS=0.137059 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=1.813e-06 SB=4.51e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=0 PANW8=3.348e-15 PANW9=2.48e-14 PANW10=3.72e-14
XMMP0 N_OUT_MMP0_d N_A_MMP0_g N_VDD_MMP0_s N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=1.8e-06 AD=7.011e-13 AS=8.136e-13 PD=2.579e-06 PS=4.504e-06 NRD=0.215556
+ NRS=0.126111 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=4.52e-07
+ SB=1.812e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=2.356e-15 PANW8=1.24e-13 PANW9=3.1744e-14 PANW10=7.44e-14
XMMP1 N_OUT_MMP0_d N_C_MMP1_g NET8 N_VDD_D0_noxref_neg PFET L=6.2e-08 W=1.8e-06
+ AD=7.011e-13 AS=4.122e-13 PD=2.579e-06 PS=2.258e-06 NRD=0.217222 NRS=0.127222
+ M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.293e-06 SB=9.71e-07 SD=0
+ PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=2.356e-15 PANW8=1.24e-14
+ PANW9=1.39744e-13 PANW10=1.896e-13
XMMP4 NET8 N_B_MMP4_g N_VDD_MMP4_s N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=1.8e-06 AD=4.122e-13 AS=8.118e-13 PD=2.258e-06 PS=4.502e-06 NRD=0.127222
+ NRS=0.125556 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.813e-06
+ SB=4.51e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=2.356e-15 PANW8=1.24e-13 PANW9=3.1744e-14 PANW10=7.44e-14
*
.include "OAI12.pex.sp.OAI12.pxi"
*
.ends
*
*
