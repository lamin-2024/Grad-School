* File: XOR2.pex.sp
* Created: Sat Nov  2 16:54:38 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.include "XOR2.pex.sp.pex"
.subckt XOR2  GND! VZ OUT VDD! VB VA
* 
* VA	VA
* VB	VB
* VDD!	VDD!
* OUT	OUT
* VZ	VZ
* GND!	GND!
XD0_noxref N_GND!_D0_noxref_pos N_VDD!_D0_noxref_neg DIODENWX  AREA=1.26612e-11
+ PERIM=1.4366e-05
XMMN1 N_VZ_MMN1_d N_VB_MMN1_g N_GND!_MMN1_s N_GND!_D0_noxref_pos NFET L=6.2e-08
+ W=1.7e-06 AD=3.825e-13 AS=7.65e-13 PD=2.15e-06 PS=4.3e-06 NRD=0.132353
+ NRS=0.132353 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=4.5e-07
+ SB=2.816e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=6.2e-17 PANW6=6.2e-15
+ PANW7=1.24e-14 PANW8=1.24e-14 PANW9=2.48e-14 PANW10=3.72e-14
XMMN0 N_VZ_MMN1_d N_VA_MMN0_g N_GND!_MMN0_s N_GND!_D0_noxref_pos NFET L=6.2e-08
+ W=1.7e-06 AD=3.825e-13 AS=3.7485e-13 PD=2.15e-06 PS=2.141e-06 NRD=0.132353
+ NRS=0.132353 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=9.62e-07
+ SB=2.304e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=6.2e-17 PANW6=6.2e-15
+ PANW7=1.24e-14 PANW8=1.24e-14 PANW9=2.48e-14 PANW10=3.72e-14
XMMN2 N_OUT_MMN2_d N_VZ_MMN2_g N_GND!_MMN0_s N_GND!_D0_noxref_pos NFET L=6.2e-08
+ W=1.7e-06 AD=3.9015e-13 AS=3.7485e-13 PD=2.159e-06 PS=2.141e-06 NRD=0.132353
+ NRS=0.127059 M=1 NF=1 CNR_SWITCH=1 PCCRIT=0 PAR=1 PTWELL=0 SA=1.465e-06
+ SB=1.801e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=6.2e-17 PANW6=6.2e-15
+ PANW7=1.24e-14 PANW8=1.24e-14 PANW9=2.48e-14 PANW10=3.72e-14
XMMN3 N_OUT_MMN2_d N_VA_MMN3_g NET25 N_GND!_D0_noxref_pos NFET L=6.2e-08
+ W=1.7e-06 AD=3.9015e-13 AS=6.528e-13 PD=2.159e-06 PS=2.468e-06 NRD=0.137647
+ NRS=0.225882 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.986e-06
+ SB=1.28e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=6.2e-17 PANW6=6.2e-15
+ PANW7=1.24e-14 PANW8=1.24e-14 PANW9=2.48e-14 PANW10=3.72e-14
XMMN4 NET25 N_VB_MMN4_g N_GND!_MMN4_s N_GND!_D0_noxref_pos NFET L=6.2e-08
+ W=1.7e-06 AD=6.528e-13 AS=7.65e-13 PD=2.468e-06 PS=4.3e-06 NRD=0.225882
+ NRS=0.132353 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=2.816e-06
+ SB=4.5e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=6.2e-17 PANW6=6.2e-15
+ PANW7=1.24e-14 PANW8=1.24e-14 PANW9=2.48e-14 PANW10=3.72e-14
XMMP0 N_VZ_MMP0_d N_VB_MMP0_g NET26 N_VDD!_D0_noxref_neg PFET L=6.2e-08
+ W=1.8e-06 AD=8.1e-13 AS=4.05e-13 PD=4.5e-06 PS=2.25e-06 NRD=0.125 NRS=0.125
+ M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=4.5e-07 SB=2.816e-06 SD=0
+ PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=1.674e-15 PANW6=6.2e-15 PANW7=1.24e-14
+ PANW8=1.34478e-13 PANW9=4.96e-14 PANW10=7.44e-14
XMMP1 NET26 N_VA_MMP1_g N_VDD!_MMP1_s N_VDD!_D0_noxref_neg PFET L=6.2e-08
+ W=1.8e-06 AD=4.05e-13 AS=3.969e-13 PD=2.25e-06 PS=2.241e-06 NRD=0.125 NRS=0.12
+ M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=9.62e-07 SB=2.304e-06 SD=0
+ PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=1.674e-15 PANW6=6.2e-15 PANW7=1.24e-14
+ PANW8=2.2878e-14 PANW9=1.486e-13 PANW10=8.7e-14
XMMP4 N_NET15_MMP4_d N_VZ_MMP4_g N_VDD!_MMP1_s N_VDD!_D0_noxref_neg PFET
+ L=6.2e-08 W=1.8e-06 AD=4.131e-13 AS=3.969e-13 PD=2.259e-06 PS=2.241e-06
+ NRD=0.125 NRS=0.125 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.465e-06
+ SB=1.801e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=1.674e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=2.2878e-14 PANW9=4.96e-14 PANW10=1.86e-13
XMMP2 N_OUT_MMP2_d N_VA_MMP2_g N_NET15_MMP4_d N_VDD!_D0_noxref_neg PFET
+ L=6.2e-08 W=1.8e-06 AD=6.912e-13 AS=4.131e-13 PD=2.568e-06 PS=2.259e-06
+ NRD=0.213333 NRS=0.13 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1
+ SA=1.986e-06 SB=1.28e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=1.674e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=2.2878e-14 PANW9=4.96e-14 PANW10=1.86e-13
XMMP3 N_OUT_MMP2_d N_VB_MMP3_g N_NET15_MMP3_s N_VDD!_D0_noxref_neg PFET
+ L=6.2e-08 W=1.8e-06 AD=6.912e-13 AS=8.1e-13 PD=2.568e-06 PS=4.5e-06
+ NRD=0.213333 NRS=0.125 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1
+ SA=2.816e-06 SB=4.5e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=1.674e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.34478e-13 PANW9=4.96e-14 PANW10=7.44e-14
c_224 NET25 0 0.00300963f
*
.include "XOR2.pex.sp.XOR2.pxi"
*
.ends
*
*
