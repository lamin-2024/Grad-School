* File: OAI22.pex.sp
* Created: Sat Nov  2 23:04:56 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.include "OAI22.pex.sp.pex"
.subckt OAI22  OUT VSS VDD VA VB VD VC
* 
* VC	VC
* VD	VD
* VB	VB
* VA	VA
* VDD	VDD
* VSS	VSS
* OUT	OUT
XD0_noxref N_VSS_D0_noxref_pos N_VDD_D0_noxref_neg DIODENWX  AREA=1.11496e-11
+ PERIM=1.3392e-05
XMMN0 N_OUT_MMN0_d N_VA_MMN0_g N_NET22_MMN0_s N_VSS_D0_noxref_pos NFET
+ L=6.2e-08 W=1.7e-06 AD=3.9015e-13 AS=7.684e-13 PD=2.159e-06 PS=4.304e-06
+ NRD=0.137647 NRS=0.133529 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=4.52e-07 SB=2.329e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=6.2e-17
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=2.48e-14 PANW10=3.72e-14
XMMN2 N_OUT_MMN0_d N_VB_MMN2_g N_NET22_MMN2_s N_VSS_D0_noxref_pos NFET
+ L=6.2e-08 W=1.7e-06 AD=3.9015e-13 AS=6.5875e-13 PD=2.159e-06 PS=2.475e-06
+ NRD=0.132353 NRS=0.338235 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=9.73e-07 SB=1.808e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=6.2e-17
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=2.48e-14 PANW10=3.72e-14
XMMN3 N_NET22_MMN2_s N_VD_MMN3_g N_VSS_MMN3_s N_VSS_D0_noxref_pos NFET
+ L=6.2e-08 W=1.7e-06 AD=6.5875e-13 AS=3.91e-13 PD=2.475e-06 PS=2.16e-06
+ NRD=0.117647 NRS=0.136471 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=1.81e-06 SB=9.71e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=6.2e-17
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=2.48e-14 PANW10=3.72e-14
XMMN1 N_NET22_MMN1_d N_VC_MMN1_g N_VSS_MMN3_s N_VSS_D0_noxref_pos NFET
+ L=6.2e-08 W=1.7e-06 AD=7.633e-13 AS=3.91e-13 PD=4.298e-06 PS=2.16e-06
+ NRD=0.131765 NRS=0.134118 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=2.332e-06 SB=4.49e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=6.2e-17
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=2.48e-14 PANW10=3.72e-14
XMMP0 NET8 N_VA_MMP0_g N_VDD_MMP0_s N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=1.8e-06 AD=4.131e-13 AS=8.136e-13 PD=2.259e-06 PS=4.504e-06 NRD=0.1275
+ NRS=0.126111 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=4.52e-07
+ SB=2.329e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=1.674e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.34478e-13 PANW9=4.96e-14 PANW10=7.44e-14
XMMP1 N_OUT_MMP1_d N_VB_MMP1_g NET8 N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=1.8e-06 AD=6.975e-13 AS=4.131e-13 PD=2.575e-06 PS=2.259e-06 NRD=0.213333
+ NRS=0.1275 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=9.73e-07
+ SB=1.808e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=1.674e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=2.2878e-14 PANW9=1.324e-13 PANW10=1.032e-13
XMMP3 N_OUT_MMP1_d N_VD_MMP3_g NET024 N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=1.8e-06 AD=6.975e-13 AS=4.14e-13 PD=2.575e-06 PS=2.26e-06 NRD=0.217222
+ NRS=0.127778 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.81e-06
+ SB=9.71e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=1.674e-15 PANW6=6.2e-15
+ PANW7=1.24e-14 PANW8=2.2878e-14 PANW9=1.594e-13 PANW10=7.62e-14
XMMP2 NET024 N_VC_MMP2_g N_VDD_MMP2_s N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=1.8e-06 AD=4.14e-13 AS=8.082e-13 PD=2.26e-06 PS=4.498e-06 NRD=0.127778
+ NRS=0.125556 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=2.332e-06
+ SB=4.49e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=1.674e-15 PANW6=6.2e-15
+ PANW7=1.24e-14 PANW8=1.34478e-13 PANW9=4.96e-14 PANW10=7.44e-14
*
.include "OAI22.pex.sp.OAI22.pxi"
*
.ends
*
*
