* File: XOR2.pex.sp
* Created: Mon Dec  2 11:45:25 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.include "XOR2.pex.sp.pex"
.subckt XOR2  VSS Z OUT VDD B A
* 
* A	A
* B	B
* VDD	VDD
* OUT	OUT
* Z	Z
* VSS	VSS
XD0_noxref N_VSS_D0_noxref_pos N_VDD_D0_noxref_neg DIODENWX  AREA=1.5785e-11
+ PERIM=1.59e-05
XMMN1 N_Z_MMN1_d N_B_MMN1_g N_VSS_MMN1_s N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=1.7e-06 AD=3.5445e-13 AS=8.636e-13 PD=2.117e-06 PS=4.416e-06 NRD=0.123529
+ NRS=0.166471 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=5.08e-07
+ SB=2.79e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=3.348e-15 PANW9=2.48e-14 PANW10=3.72e-14
XMMN0 N_Z_MMN1_d N_A_MMN0_g N_VSS_MMN0_s N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=1.7e-06 AD=3.5445e-13 AS=3.7485e-13 PD=2.117e-06 PS=2.141e-06 NRD=0.121765
+ NRS=0.132353 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=9.87e-07
+ SB=2.311e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=3.348e-15 PANW9=2.48e-14 PANW10=3.72e-14
XMMN2 N_OUT_MMN2_d N_Z_MMN2_g N_VSS_MMN0_s N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=1.7e-06 AD=3.893e-13 AS=3.7485e-13 PD=2.158e-06 PS=2.141e-06 NRD=0.131765
+ NRS=0.127059 M=1 NF=1 CNR_SWITCH=1 PCCRIT=0 PAR=1 PTWELL=0 SA=1.49e-06
+ SB=1.808e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=3.348e-15 PANW9=2.48e-14 PANW10=3.72e-14
XMMN3 N_OUT_MMN2_d N_A_MMN3_g NET25 N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=1.7e-06 AD=3.893e-13 AS=6.596e-13 PD=2.158e-06 PS=2.476e-06 NRD=0.137647
+ NRS=0.228235 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=2.01e-06
+ SB=1.288e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=3.348e-15 PANW9=2.48e-14 PANW10=3.72e-14
XMMN4 NET25 N_B_MMN4_g N_VSS_MMN4_s N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=1.7e-06 AD=6.596e-13 AS=7.65e-13 PD=2.476e-06 PS=4.3e-06 NRD=0.228235
+ NRS=0.132353 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=2.848e-06
+ SB=4.5e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=3.348e-15 PANW9=2.48e-14 PANW10=3.72e-14
XMMP0 N_Z_MMP0_d N_B_MMP0_g NET26 N_VDD_D0_noxref_neg PFET L=6.2e-08 W=1.8e-06
+ AD=9.144e-13 AS=3.753e-13 PD=4.616e-06 PS=2.217e-06 NRD=0.157222 NRS=0.115833
+ M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=5.08e-07 SB=2.79e-06 SD=0
+ PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=2.356e-15 PANW8=1.24e-13
+ PANW9=3.1744e-14 PANW10=7.44e-14
XMMP1 NET26 N_A_MMP1_g N_VDD_MMP1_s N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=1.8e-06 AD=3.753e-13 AS=3.969e-13 PD=2.217e-06 PS=2.241e-06 NRD=0.115833
+ NRS=0.12 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=9.87e-07
+ SB=2.311e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=2.356e-15 PANW8=1.24e-14 PANW9=1.09144e-13 PANW10=1.086e-13
XMMP4 N_NET15_MMP4_d N_Z_MMP4_g N_VDD_MMP1_s N_VDD_D0_noxref_neg PFET
+ L=6.2e-08 W=1.8e-06 AD=4.122e-13 AS=3.969e-13 PD=2.258e-06 PS=2.241e-06
+ NRD=0.124444 NRS=0.125 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1
+ SA=1.49e-06 SB=1.808e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=2.356e-15 PANW8=1.24e-14 PANW9=3.1744e-14 PANW10=1.86e-13
XMMP2 N_OUT_MMP2_d N_A_MMP2_g N_NET15_MMP4_d N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=1.8e-06 AD=6.984e-13 AS=4.122e-13 PD=2.576e-06 PS=2.258e-06 NRD=0.213889
+ NRS=0.13 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=2.01e-06
+ SB=1.288e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=2.356e-15 PANW8=1.24e-14 PANW9=3.1744e-14 PANW10=1.86e-13
XMMP3 N_OUT_MMP2_d N_B_MMP3_g N_NET15_MMP3_s N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=1.8e-06 AD=6.984e-13 AS=8.1e-13 PD=2.576e-06 PS=4.5e-06 NRD=0.217222
+ NRS=0.125 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=2.848e-06
+ SB=4.5e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=2.356e-15 PANW8=1.24e-13 PANW9=3.1744e-14 PANW10=7.44e-14
*
.include "XOR2.pex.sp.XOR2.pxi"
*
.ends
*
*
